module PacifikerClaws(
  input CLK,
  output RST,
  output SCL,
  output DC,
  output MOSI,
  output CS
 );

 // LCD Command names from Pulse View
 localparam SLPOUT  = 8'h11;
 localparam FRMCTR1 = 8'hB1;
 localparam FRMCTR2 = 8'hB2;
 localparam FRMCTR3 = 8'hB3;
 localparam INVCTR  = 8'hB4;
 localparam PWCTR1  = 8'hC0;
 localparam PWCTR2  = 8'hC1;
 localparam PWCTR3  = 8'hC2;
 localparam PWCTR4  = 8'hC3;
 localparam PWCTR5  = 8'hC4;
 localparam VMCTR1  = 8'hC5;
 localparam GMCTRP1 = 8'hE0;
 localparam GMCTRN1 = 8'hE1;
 localparam PWCTR6  = 8'hFC;
 localparam COLMOD  = 8'h3A;
 localparam MADCTL  = 8'h36;
 localparam INVON   = 8'h21;
 localparam DISPON  = 8'h29;
 localparam CASET   = 8'h2A;
 localparam RASET   = 8'h2B;
 localparam RAMWR   = 8'h2C;

 localparam init = 6'd0;
 localparam actRst = 6'd1;
 localparam drst = 6'd2;
 localparam ddrst = 6'd3;
 localparam lc = 6'd4;
 localparam ldc = 6'd5;
 localparam sm = 6'd6;
 localparam lcs = 6'd7;
 localparam slb = 6'd8;
 localparam rcs = 6'd9;
 localparam send = 6'd10;
 localparam rdc = 6'd11;
 localparam lp = 6'd12;
 localparam dsleep = 6'd13;
 localparam dpcmd = 6'd14;
 localparam dmw_c = 6'd15;
 localparam dmw_p = 6'd16;
 localparam dcrg_p = 6'd17;
 localparam dfrmctr3_c = 6'd18;
 localparam dfrmctr3_p = 6'd19;
 localparam dgmctr_c = 6'd20;
 localparam dgmctr_p = 6'd21;
 localparam dcr_c = 6'd22;
 localparam dcr_p = 6'd23;

 localparam actRst_d = 16'd23817;
 localparam dactRst_d = 16'd20858;
 localparam sleep = 16'd20848;
 localparam pcmd = 12'd36; // 3us post cmd delay
 localparam mw_c = 12'd480; // 40us post memory write
 localparam mw_p = 12'd72; // memory write param
 localparam crg = 12'd36; //CASET/RASET/Gamma+/- del.
 localparam frmctr3 = 12'd36;
 localparam gmctr = 12'd36; // 3us for gamma ctr
 localparam cr = 12'd36; // 3us for caset raset

 reg rst, scl, dc, mosi, cs;
 reg [5:0] state;
 reg [15:0] delay;

 reg [7:0] data;
 reg [2:0] bit_counter; 
 
 reg [15:0] pixel_data;
 reg [3:0] pixel_bit_counter;

 reg [7:0] cmd [0:21];
 reg [4:0] cmd_counter;

 reg [7:0] params [0:67];
 reg [6:0] param_counter;

 reg [13:0] params_left;

 reg [7:0] picture_data [0:7599];
 reg [12:0] pic_pointer;

 initial
 begin
  state = 6'd0;
  scl = 1'b1;

  cmd[0]  = SLPOUT;
  cmd[1]  = FRMCTR1;
  cmd[2]  = FRMCTR2;
  cmd[3]  = FRMCTR3;
  cmd[4]  = INVCTR;
  cmd[5]  = PWCTR1;
  cmd[6]  = PWCTR2;
  cmd[7]  = PWCTR3;
  cmd[8]  = PWCTR4;
  cmd[9]  = PWCTR5;
  cmd[10] = VMCTR1;
  cmd[11] = GMCTRP1;
  cmd[12] = GMCTRN1;
  cmd[13] = PWCTR6;
  cmd[14] = COLMOD;
  cmd[15] = MADCTL;
  cmd[16] = INVON;
  cmd[17] = DISPON;
  cmd[18] = CASET;
  cmd[19] = RASET;
  cmd[20] = RAMWR; 
  cmd[21] = 8'h00; //NOP
  cmd_counter = 5'b0;

  params[0]  = 8'h05;
  params[1]  = 8'h3C;
  params[2]  = 8'h3C;
  params[3]  = 8'h05;
  params[4]  = 8'h3C;
  params[5]  = 8'h3C;
  params[6]  = 8'h05;
  params[7]  = 8'h3C;
  params[8]  = 8'h3C;
  params[9]  = 8'h05;
  params[10] = 8'h3C;
  params[11] = 8'h3C;
  params[12] = 8'h03;
  params[13] = 8'hAB;
  params[14] = 8'h0B;
  params[15] = 8'h04;
  params[16] = 8'hC5;
  params[17] = 8'h0D;
  params[18] = 8'h00;
  params[19] = 8'h8D;
  params[20] = 8'h6A;
  params[21] = 8'h8D;
  params[22] = 8'hEE;
  params[23] = 8'h0F;
  params[24] = 8'h07;
  params[25] = 8'h0E;
  params[26] = 8'h08;
  params[27] = 8'h07;
  params[28] = 8'h10;
  params[29] = 8'h07;
  params[30] = 8'h02;
  params[31] = 8'h07;
  params[32] = 8'h09;
  params[33] = 8'h0F;
  params[34] = 8'h25;
  params[35] = 8'h36;
  params[36] = 8'h00;
  params[37] = 8'h08;
  params[38] = 8'h04;
  params[39] = 8'h10;
  params[40] = 8'h0A;
  params[41] = 8'h0D;
  params[42] = 8'h08;
  params[43] = 8'h07;
  params[44] = 8'h0F;
  params[45] = 8'h07;
  params[46] = 8'h02;
  params[47] = 8'h07;
  params[48] = 8'h09;
  params[49] = 8'h0F;
  params[50] = 8'h25;
  params[51] = 8'h35;
  params[52] = 8'h00;
  params[53] = 8'h09;
  params[54] = 8'h04;
  params[55] = 8'h10;
  params[56] = 8'h80;
  params[57] = 8'h05;
  params[58] = 8'h78;
  params[59] = 8'h00;
  params[60] = 8'h2B;
  params[61] = 8'h00;
  params[62] = 8'h76;// 002B - 0076
  params[63] = 8'h00;
  params[64] = 8'h29;
  params[65] = 8'h00;
  params[66] = 8'h5A;// 0029 - 005A
  //params[67] = 8'hC7;// Limish Color

  param_counter = 7'b00;
  params_left = 14'd0;

  data = 8'h00;
  bit_counter = 3'b111;

  pixel_data = 16'h00_00;
  pixel_bit_counter = 4'b1111;

  picture_data[ 0 ] = 8'hCD;   
  picture_data[ 1 ] = 8'hF7;
  picture_data[ 2 ] = 8'h39;
  picture_data[ 3 ] = 8'hA6;
  picture_data[ 4 ] = 8'h18;
  picture_data[ 5 ] = 8'hC2;
  picture_data[ 6 ] = 8'h29;
  picture_data[ 7 ] = 8'h64;
  picture_data[ 8 ] = 8'h19;
  picture_data[ 9 ] = 8'h02;
  picture_data[ 10 ] = 8'h19;
  picture_data[ 11 ] = 8'h22;
  picture_data[ 12 ] = 8'h18;
  picture_data[ 13 ] = 8'hE1;
  picture_data[ 14 ] = 8'h41;
  picture_data[ 15 ] = 8'hC4;
  picture_data[ 16 ] = 8'h7B;
  picture_data[ 17 ] = 8'h49;
  picture_data[ 18 ] = 8'hA4;
  picture_data[ 19 ] = 8'hAE;
  picture_data[ 20 ] = 8'hD6;
  picture_data[ 21 ] = 8'h74;
  picture_data[ 22 ] = 8'hEF;
  picture_data[ 23 ] = 8'h37;
  picture_data[ 24 ] = 8'h5A;
  picture_data[ 25 ] = 8'hC6;
  picture_data[ 26 ] = 8'h9C;
  picture_data[ 27 ] = 8'hEE;
  picture_data[ 28 ] = 8'hD6;
  picture_data[ 29 ] = 8'h75;
  picture_data[ 30 ] = 8'h8C;
  picture_data[ 31 ] = 8'h2C;
  picture_data[ 32 ] = 8'h7B;
  picture_data[ 33 ] = 8'h6B;
  picture_data[ 34 ] = 8'h73;
  picture_data[ 35 ] = 8'h09;
  picture_data[ 36 ] = 8'hCD;
  picture_data[ 37 ] = 8'h93;
  picture_data[ 38 ] = 8'hB4;
  picture_data[ 39 ] = 8'hF0;
  picture_data[ 40 ] = 8'hAC;
  picture_data[ 41 ] = 8'hF0;
  picture_data[ 42 ] = 8'hD6;
  picture_data[ 43 ] = 8'h96;
  picture_data[ 44 ] = 8'hB5;
  picture_data[ 45 ] = 8'hD4;
  picture_data[ 46 ] = 8'hAD;
  picture_data[ 47 ] = 8'hB4;
  picture_data[ 48 ] = 8'h84;
  picture_data[ 49 ] = 8'h4F;
  picture_data[ 50 ] = 8'h73;
  picture_data[ 51 ] = 8'h8B;
  picture_data[ 52 ] = 8'h63;
  picture_data[ 53 ] = 8'h29;
  picture_data[ 54 ] = 8'h94;
  picture_data[ 55 ] = 8'hAF;
  picture_data[ 56 ] = 8'h94;
  picture_data[ 57 ] = 8'hAF;
  picture_data[ 58 ] = 8'hCE;
  picture_data[ 59 ] = 8'h56;
  picture_data[ 60 ] = 8'h9C;
  picture_data[ 61 ] = 8'hD1;
  picture_data[ 62 ] = 8'h39;
  picture_data[ 63 ] = 8'hA5;
  picture_data[ 64 ] = 8'h39;
  picture_data[ 65 ] = 8'h64;
  picture_data[ 66 ] = 8'h20;
  picture_data[ 67 ] = 8'hE2;
  picture_data[ 68 ] = 8'h31;
  picture_data[ 69 ] = 8'hA5;
  picture_data[ 70 ] = 8'h21;
  picture_data[ 71 ] = 8'h43;
  picture_data[ 72 ] = 8'h39;
  picture_data[ 73 ] = 8'hE5;
  picture_data[ 74 ] = 8'h6B;
  picture_data[ 75 ] = 8'h4B;
  picture_data[ 76 ] = 8'h39;
  picture_data[ 77 ] = 8'h23;
  picture_data[ 78 ] = 8'h28;
  picture_data[ 79 ] = 8'hC3;
  picture_data[ 80 ] = 8'h10;
  picture_data[ 81 ] = 8'h62;
  picture_data[ 82 ] = 8'h10;
  picture_data[ 83 ] = 8'hA3;
  picture_data[ 84 ] = 8'h08;
  picture_data[ 85 ] = 8'h82;
  picture_data[ 86 ] = 8'h08;
  picture_data[ 87 ] = 8'hC2;
  picture_data[ 88 ] = 8'h09;
  picture_data[ 89 ] = 8'h04;
  picture_data[ 90 ] = 8'h01;
  picture_data[ 91 ] = 8'hC6;
  picture_data[ 92 ] = 8'h0A;
  picture_data[ 93 ] = 8'hA9;
  picture_data[ 94 ] = 8'h1B;
  picture_data[ 95 ] = 8'hAD;
  picture_data[ 96 ] = 8'h02;
  picture_data[ 97 ] = 8'hA9;
  picture_data[ 98 ] = 8'h02;
  picture_data[ 99 ] = 8'hAA;
  picture_data[ 100 ] = 8'h01;
  picture_data[ 101 ] = 8'hE7;
  picture_data[ 102 ] = 8'h09;
  picture_data[ 103 ] = 8'hA6;
  picture_data[ 104 ] = 8'h3A;
  picture_data[ 105 ] = 8'hA8;
  picture_data[ 106 ] = 8'h3A;
  picture_data[ 107 ] = 8'h47;
  picture_data[ 108 ] = 8'h39;
  picture_data[ 109 ] = 8'hC7;
  picture_data[ 110 ] = 8'h18;
  picture_data[ 111 ] = 8'hE4;
  picture_data[ 112 ] = 8'h19;
  picture_data[ 113 ] = 8'h03;
  picture_data[ 114 ] = 8'h10;
  picture_data[ 115 ] = 8'hC2;
  picture_data[ 116 ] = 8'h21;
  picture_data[ 117 ] = 8'h03;
  picture_data[ 118 ] = 8'h31;
  picture_data[ 119 ] = 8'h44;
  picture_data[ 120 ] = 8'h29;
  picture_data[ 121 ] = 8'h22;
  picture_data[ 122 ] = 8'h20;
  picture_data[ 123 ] = 8'hE1;
  picture_data[ 124 ] = 8'h41;
  picture_data[ 125 ] = 8'hE6;
  picture_data[ 126 ] = 8'h41;
  picture_data[ 127 ] = 8'hA6;
  picture_data[ 128 ] = 8'h41;
  picture_data[ 129 ] = 8'hC5;
  picture_data[ 130 ] = 8'h4A;
  picture_data[ 131 ] = 8'h06;
  picture_data[ 132 ] = 8'h5A;
  picture_data[ 133 ] = 8'hA8;
  picture_data[ 134 ] = 8'h5A;
  picture_data[ 135 ] = 8'hC8;
  picture_data[ 136 ] = 8'h20;
  picture_data[ 137 ] = 8'hE1;
  picture_data[ 138 ] = 8'h4A;
  picture_data[ 139 ] = 8'h25;
  picture_data[ 140 ] = 8'h4A;
  picture_data[ 141 ] = 8'h05;
  picture_data[ 142 ] = 8'h21;
  picture_data[ 143 ] = 8'h00;
  picture_data[ 144 ] = 8'h29;
  picture_data[ 145 ] = 8'h00;
  picture_data[ 146 ] = 8'h41;
  picture_data[ 147 ] = 8'h82;
  picture_data[ 148 ] = 8'h52;
  picture_data[ 149 ] = 8'h04;
  picture_data[ 150 ] = 8'h7B;
  picture_data[ 151 ] = 8'h6A;
  picture_data[ 152 ] = 8'hBD;
  picture_data[ 153 ] = 8'h95;
  picture_data[ 154 ] = 8'h62;
  picture_data[ 155 ] = 8'hCA;
  picture_data[ 156 ] = 8'h29;
  picture_data[ 157 ] = 8'h44;
  picture_data[ 158 ] = 8'h19;
  picture_data[ 159 ] = 8'h23;
  picture_data[ 160 ] = 8'h21;
  picture_data[ 161 ] = 8'h43;
  picture_data[ 162 ] = 8'h29;
  picture_data[ 163 ] = 8'h64;
  picture_data[ 164 ] = 8'h29;
  picture_data[ 165 ] = 8'h63;
  picture_data[ 166 ] = 8'h29;
  picture_data[ 167 ] = 8'h42;
  picture_data[ 168 ] = 8'hBD;
  picture_data[ 169 ] = 8'h92;
  picture_data[ 170 ] = 8'hDE;
  picture_data[ 171 ] = 8'h96;
  picture_data[ 172 ] = 8'hBD;
  picture_data[ 173 ] = 8'hB2;
  picture_data[ 174 ] = 8'hD6;
  picture_data[ 175 ] = 8'h54;
  picture_data[ 176 ] = 8'h42;
  picture_data[ 177 ] = 8'h03;
  picture_data[ 178 ] = 8'h63;
  picture_data[ 179 ] = 8'h07;
  picture_data[ 180 ] = 8'hB5;
  picture_data[ 181 ] = 8'h92;
  picture_data[ 182 ] = 8'h52;
  picture_data[ 183 ] = 8'h66;
  picture_data[ 184 ] = 8'h42;
  picture_data[ 185 ] = 8'h05;
  picture_data[ 186 ] = 8'h73;
  picture_data[ 187 ] = 8'h4A;
  picture_data[ 188 ] = 8'h94;
  picture_data[ 189 ] = 8'h0D;
  picture_data[ 190 ] = 8'h8B;
  picture_data[ 191 ] = 8'hAB;
  picture_data[ 192 ] = 8'h94;
  picture_data[ 193 ] = 8'h4D;
  picture_data[ 194 ] = 8'h8C;
  picture_data[ 195 ] = 8'h2D;
  picture_data[ 196 ] = 8'h52;
  picture_data[ 197 ] = 8'hA8;
  picture_data[ 198 ] = 8'h52;
  picture_data[ 199 ] = 8'hE9;
  picture_data[ 200 ] = 8'h4A;
  picture_data[ 201 ] = 8'hA8;
  picture_data[ 202 ] = 8'h52;
  picture_data[ 203 ] = 8'hA8;
  picture_data[ 204 ] = 8'h5A;
  picture_data[ 205 ] = 8'hE9;
  picture_data[ 206 ] = 8'h52;
  picture_data[ 207 ] = 8'h87;
  picture_data[ 208 ] = 8'h5A;
  picture_data[ 209 ] = 8'hC8;
  picture_data[ 210 ] = 8'h7B;
  picture_data[ 211 ] = 8'hCC;
  picture_data[ 212 ] = 8'h31;
  picture_data[ 213 ] = 8'h84;
  picture_data[ 214 ] = 8'h29;
  picture_data[ 215 ] = 8'h43;
  picture_data[ 216 ] = 8'h41;
  picture_data[ 217 ] = 8'hC5;
  picture_data[ 218 ] = 8'h52;
  picture_data[ 219 ] = 8'h68;
  picture_data[ 220 ] = 8'h31;
  picture_data[ 221 ] = 8'hC5;
  picture_data[ 222 ] = 8'h21;
  picture_data[ 223 ] = 8'h23;
  picture_data[ 224 ] = 8'h29;
  picture_data[ 225 ] = 8'h43;
  picture_data[ 226 ] = 8'h29;
  picture_data[ 227 ] = 8'h02;
  picture_data[ 228 ] = 8'h39;
  picture_data[ 229 ] = 8'h44;
  picture_data[ 230 ] = 8'h28;
  picture_data[ 231 ] = 8'hC2;
  picture_data[ 232 ] = 8'h10;
  picture_data[ 233 ] = 8'h42;
  picture_data[ 234 ] = 8'h10;
  picture_data[ 235 ] = 8'h83;
  picture_data[ 236 ] = 8'h18;
  picture_data[ 237 ] = 8'hE3;
  picture_data[ 238 ] = 8'h19;
  picture_data[ 239 ] = 8'h44;
  picture_data[ 240 ] = 8'h01;
  picture_data[ 241 ] = 8'h45;
  picture_data[ 242 ] = 8'h02;
  picture_data[ 243 ] = 8'h08;
  picture_data[ 244 ] = 8'h03;
  picture_data[ 245 ] = 8'h0B;
  picture_data[ 246 ] = 8'h35;
  picture_data[ 247 ] = 8'h53;
  picture_data[ 248 ] = 8'h2C;
  picture_data[ 249 ] = 8'hB2;
  picture_data[ 250 ] = 8'h0B;
  picture_data[ 251 ] = 8'h4C;
  picture_data[ 252 ] = 8'h0A;
  picture_data[ 253 ] = 8'h28;
  picture_data[ 254 ] = 8'h1A;
  picture_data[ 255 ] = 8'h07;
  picture_data[ 256 ] = 8'h19;
  picture_data[ 257 ] = 8'hC5;
  picture_data[ 258 ] = 8'h19;
  picture_data[ 259 ] = 8'h64;
  picture_data[ 260 ] = 8'h21;
  picture_data[ 261 ] = 8'h45;
  picture_data[ 262 ] = 8'h18;
  picture_data[ 263 ] = 8'hC3;
  picture_data[ 264 ] = 8'h19;
  picture_data[ 265 ] = 8'h03;
  picture_data[ 266 ] = 8'h19;
  picture_data[ 267 ] = 8'h23;
  picture_data[ 268 ] = 8'h18;
  picture_data[ 269 ] = 8'hC2;
  picture_data[ 270 ] = 8'h29;
  picture_data[ 271 ] = 8'h23;
  picture_data[ 272 ] = 8'h31;
  picture_data[ 273 ] = 8'hA4;
  picture_data[ 274 ] = 8'h29;
  picture_data[ 275 ] = 8'h63;
  picture_data[ 276 ] = 8'h21;
  picture_data[ 277 ] = 8'h02;
  picture_data[ 278 ] = 8'h20;
  picture_data[ 279 ] = 8'hE2;
  picture_data[ 280 ] = 8'h18;
  picture_data[ 281 ] = 8'hC1;
  picture_data[ 282 ] = 8'h41;
  picture_data[ 283 ] = 8'hE5;
  picture_data[ 284 ] = 8'h42;
  picture_data[ 285 ] = 8'h06;
  picture_data[ 286 ] = 8'h29;
  picture_data[ 287 ] = 8'h42;
  picture_data[ 288 ] = 8'h31;
  picture_data[ 289 ] = 8'h63;
  picture_data[ 290 ] = 8'h52;
  picture_data[ 291 ] = 8'h46;
  picture_data[ 292 ] = 8'h29;
  picture_data[ 293 ] = 8'h21;
  picture_data[ 294 ] = 8'h52;
  picture_data[ 295 ] = 8'h25;
  picture_data[ 296 ] = 8'h73;
  picture_data[ 297 ] = 8'h49;
  picture_data[ 298 ] = 8'hBD;
  picture_data[ 299 ] = 8'h51;
  picture_data[ 300 ] = 8'hD6;
  picture_data[ 301 ] = 8'h14;
  picture_data[ 302 ] = 8'hCD;
  picture_data[ 303 ] = 8'hD3;
  picture_data[ 304 ] = 8'hB5;
  picture_data[ 305 ] = 8'h53;
  picture_data[ 306 ] = 8'h63;
  picture_data[ 307 ] = 8'h0A;
  picture_data[ 308 ] = 8'h10;
  picture_data[ 309 ] = 8'hA1;
  picture_data[ 310 ] = 8'h21;
  picture_data[ 311 ] = 8'h43;
  picture_data[ 312 ] = 8'h29;
  picture_data[ 313 ] = 8'hC5;
  picture_data[ 314 ] = 8'h19;
  picture_data[ 315 ] = 8'h02;
  picture_data[ 316 ] = 8'h29;
  picture_data[ 317 ] = 8'h63;
  picture_data[ 318 ] = 8'h21;
  picture_data[ 319 ] = 8'h22;
  picture_data[ 320 ] = 8'h52;
  picture_data[ 321 ] = 8'h66;
  picture_data[ 322 ] = 8'hAD;
  picture_data[ 323 ] = 8'h31;
  picture_data[ 324 ] = 8'hCE;
  picture_data[ 325 ] = 8'h14;
  picture_data[ 326 ] = 8'hA4;
  picture_data[ 327 ] = 8'hF0;
  picture_data[ 328 ] = 8'h31;
  picture_data[ 329 ] = 8'h62;
  picture_data[ 330 ] = 8'h31;
  picture_data[ 331 ] = 8'h42;
  picture_data[ 332 ] = 8'h31;
  picture_data[ 333 ] = 8'h63;
  picture_data[ 334 ] = 8'h31;
  picture_data[ 335 ] = 8'h63;
  picture_data[ 336 ] = 8'h31;
  picture_data[ 337 ] = 8'hA4;
  picture_data[ 338 ] = 8'h4A;
  picture_data[ 339 ] = 8'h26;
  picture_data[ 340 ] = 8'h62;
  picture_data[ 341 ] = 8'hA8;
  picture_data[ 342 ] = 8'h62;
  picture_data[ 343 ] = 8'h88;
  picture_data[ 344 ] = 8'h52;
  picture_data[ 345 ] = 8'h46;
  picture_data[ 346 ] = 8'h4A;
  picture_data[ 347 ] = 8'h67;
  picture_data[ 348 ] = 8'h52;
  picture_data[ 349 ] = 8'hC9;
  picture_data[ 350 ] = 8'h3A;
  picture_data[ 351 ] = 8'h27;
  picture_data[ 352 ] = 8'h4A;
  picture_data[ 353 ] = 8'hA9;
  picture_data[ 354 ] = 8'h42;
  picture_data[ 355 ] = 8'h47;
  picture_data[ 356 ] = 8'h39;
  picture_data[ 357 ] = 8'hE5;
  picture_data[ 358 ] = 8'h5A;
  picture_data[ 359 ] = 8'hE9;
  picture_data[ 360 ] = 8'h4A;
  picture_data[ 361 ] = 8'h87;
  picture_data[ 362 ] = 8'h29;
  picture_data[ 363 ] = 8'h63;
  picture_data[ 364 ] = 8'h39;
  picture_data[ 365 ] = 8'hC5;
  picture_data[ 366 ] = 8'h39;
  picture_data[ 367 ] = 8'hC5;
  picture_data[ 368 ] = 8'h52;
  picture_data[ 369 ] = 8'hC9;
  picture_data[ 370 ] = 8'h52;
  picture_data[ 371 ] = 8'hC9;
  picture_data[ 372 ] = 8'h31;
  picture_data[ 373 ] = 8'hA4;
  picture_data[ 374 ] = 8'h29;
  picture_data[ 375 ] = 8'h42;
  picture_data[ 376 ] = 8'h29;
  picture_data[ 377 ] = 8'h02;
  picture_data[ 378 ] = 8'h31;
  picture_data[ 379 ] = 8'h23;
  picture_data[ 380 ] = 8'h10;
  picture_data[ 381 ] = 8'h60;
  picture_data[ 382 ] = 8'h18;
  picture_data[ 383 ] = 8'h81;
  picture_data[ 384 ] = 8'h18;
  picture_data[ 385 ] = 8'hA3;
  picture_data[ 386 ] = 8'h18;
  picture_data[ 387 ] = 8'hA3;
  picture_data[ 388 ] = 8'h10;
  picture_data[ 389 ] = 8'hE3;
  picture_data[ 390 ] = 8'h09;
  picture_data[ 391 ] = 8'h03;
  picture_data[ 392 ] = 8'h01;
  picture_data[ 393 ] = 8'h66;
  picture_data[ 394 ] = 8'h24;
  picture_data[ 395 ] = 8'h10;
  picture_data[ 396 ] = 8'h2E;
  picture_data[ 397 ] = 8'h99;
  picture_data[ 398 ] = 8'h3F;
  picture_data[ 399 ] = 8'h9D;
  picture_data[ 400 ] = 8'h7F;
  picture_data[ 401 ] = 8'hFF;
  picture_data[ 402 ] = 8'h24;
  picture_data[ 403 ] = 8'h51;
  picture_data[ 404 ] = 8'h02;
  picture_data[ 405 ] = 8'h28;
  picture_data[ 406 ] = 8'h11;
  picture_data[ 407 ] = 8'hE7;
  picture_data[ 408 ] = 8'h09;
  picture_data[ 409 ] = 8'h64;
  picture_data[ 410 ] = 8'h11;
  picture_data[ 411 ] = 8'h23;
  picture_data[ 412 ] = 8'h10;
  picture_data[ 413 ] = 8'hE4;
  picture_data[ 414 ] = 8'h18;
  picture_data[ 415 ] = 8'hE4;
  picture_data[ 416 ] = 8'h19;
  picture_data[ 417 ] = 8'h02;
  picture_data[ 418 ] = 8'h21;
  picture_data[ 419 ] = 8'h22;
  picture_data[ 420 ] = 8'h21;
  picture_data[ 421 ] = 8'h23;
  picture_data[ 422 ] = 8'h29;
  picture_data[ 423 ] = 8'h63;
  picture_data[ 424 ] = 8'h21;
  picture_data[ 425 ] = 8'h83;
  picture_data[ 426 ] = 8'h21;
  picture_data[ 427 ] = 8'hA3;
  picture_data[ 428 ] = 8'h29;
  picture_data[ 429 ] = 8'h84;
  picture_data[ 430 ] = 8'h39;
  picture_data[ 431 ] = 8'hC5;
  picture_data[ 432 ] = 8'h29;
  picture_data[ 433 ] = 8'h84;
  picture_data[ 434 ] = 8'h21;
  picture_data[ 435 ] = 8'h23;
  picture_data[ 436 ] = 8'h29;
  picture_data[ 437 ] = 8'h43;
  picture_data[ 438 ] = 8'h31;
  picture_data[ 439 ] = 8'h84;
  picture_data[ 440 ] = 8'h6B;
  picture_data[ 441 ] = 8'h0A;
  picture_data[ 442 ] = 8'h73;
  picture_data[ 443 ] = 8'h4A;
  picture_data[ 444 ] = 8'h5A;
  picture_data[ 445 ] = 8'h46;
  picture_data[ 446 ] = 8'h9C;
  picture_data[ 447 ] = 8'h6E;
  picture_data[ 448 ] = 8'hAC;
  picture_data[ 449 ] = 8'hCF;
  picture_data[ 450 ] = 8'hAC;
  picture_data[ 451 ] = 8'hCF;
  picture_data[ 452 ] = 8'hB5;
  picture_data[ 453 ] = 8'h30;
  picture_data[ 454 ] = 8'hCD;
  picture_data[ 455 ] = 8'hD2;
  picture_data[ 456 ] = 8'h8C;
  picture_data[ 457 ] = 8'h4F;
  picture_data[ 458 ] = 8'h4A;
  picture_data[ 459 ] = 8'h67;
  picture_data[ 460 ] = 8'h10;
  picture_data[ 461 ] = 8'hE1;
  picture_data[ 462 ] = 8'h10;
  picture_data[ 463 ] = 8'hC1;
  picture_data[ 464 ] = 8'h31;
  picture_data[ 465 ] = 8'hE5;
  picture_data[ 466 ] = 8'h42;
  picture_data[ 467 ] = 8'h47;
  picture_data[ 468 ] = 8'h21;
  picture_data[ 469 ] = 8'h43;
  picture_data[ 470 ] = 8'h18;
  picture_data[ 471 ] = 8'hC1;
  picture_data[ 472 ] = 8'h4A;
  picture_data[ 473 ] = 8'h46;
  picture_data[ 474 ] = 8'h4A;
  picture_data[ 475 ] = 8'h46;
  picture_data[ 476 ] = 8'h94;
  picture_data[ 477 ] = 8'h8F;
  picture_data[ 478 ] = 8'h9C;
  picture_data[ 479 ] = 8'hB0;
  picture_data[ 480 ] = 8'h31;
  picture_data[ 481 ] = 8'h63;
  picture_data[ 482 ] = 8'h31;
  picture_data[ 483 ] = 8'h64;
  picture_data[ 484 ] = 8'h31;
  picture_data[ 485 ] = 8'h84;
  picture_data[ 486 ] = 8'h31;
  picture_data[ 487 ] = 8'hA5;
  picture_data[ 488 ] = 8'h42;
  picture_data[ 489 ] = 8'h06;
  picture_data[ 490 ] = 8'h4A;
  picture_data[ 491 ] = 8'h47;
  picture_data[ 492 ] = 8'h4A;
  picture_data[ 493 ] = 8'h26;
  picture_data[ 494 ] = 8'h41;
  picture_data[ 495 ] = 8'hC5;
  picture_data[ 496 ] = 8'h39;
  picture_data[ 497 ] = 8'hC5;
  picture_data[ 498 ] = 8'h42;
  picture_data[ 499 ] = 8'h47;
  picture_data[ 500 ] = 8'h31;
  picture_data[ 501 ] = 8'hE6;
  picture_data[ 502 ] = 8'h29;
  picture_data[ 503 ] = 8'hC5;
  picture_data[ 504 ] = 8'h4A;
  picture_data[ 505 ] = 8'hA9;
  picture_data[ 506 ] = 8'h31;
  picture_data[ 507 ] = 8'hC5;
  picture_data[ 508 ] = 8'h29;
  picture_data[ 509 ] = 8'hA4;
  picture_data[ 510 ] = 8'h29;
  picture_data[ 511 ] = 8'hA4;
  picture_data[ 512 ] = 8'h29;
  picture_data[ 513 ] = 8'hA4;
  picture_data[ 514 ] = 8'h39;
  picture_data[ 515 ] = 8'hE5;
  picture_data[ 516 ] = 8'h42;
  picture_data[ 517 ] = 8'h27;
  picture_data[ 518 ] = 8'h39;
  picture_data[ 519 ] = 8'hC6;
  picture_data[ 520 ] = 8'h19;
  picture_data[ 521 ] = 8'h02;
  picture_data[ 522 ] = 8'h21;
  picture_data[ 523 ] = 8'h43;
  picture_data[ 524 ] = 8'h29;
  picture_data[ 525 ] = 8'h42;
  picture_data[ 526 ] = 8'h31;
  picture_data[ 527 ] = 8'h43;
  picture_data[ 528 ] = 8'h31;
  picture_data[ 529 ] = 8'h44;
  picture_data[ 530 ] = 8'h28;
  picture_data[ 531 ] = 8'hE2;
  picture_data[ 532 ] = 8'h20;
  picture_data[ 533 ] = 8'hA1;
  picture_data[ 534 ] = 8'h28;
  picture_data[ 535 ] = 8'hE2;
  picture_data[ 536 ] = 8'h20;
  picture_data[ 537 ] = 8'hE3;
  picture_data[ 538 ] = 8'h18;
  picture_data[ 539 ] = 8'hC3;
  picture_data[ 540 ] = 8'h11;
  picture_data[ 541 ] = 8'h04;
  picture_data[ 542 ] = 8'h09;
  picture_data[ 543 ] = 8'h45;
  picture_data[ 544 ] = 8'h01;
  picture_data[ 545 ] = 8'hC7;
  picture_data[ 546 ] = 8'h13;
  picture_data[ 547 ] = 8'hEF;
  picture_data[ 548 ] = 8'h3F;
  picture_data[ 549 ] = 8'h5C;
  picture_data[ 550 ] = 8'h37;
  picture_data[ 551 ] = 8'h7D;
  picture_data[ 552 ] = 8'h6F;
  picture_data[ 553 ] = 8'h9E;
  picture_data[ 554 ] = 8'h2C;
  picture_data[ 555 ] = 8'h92;
  picture_data[ 556 ] = 8'h01;
  picture_data[ 557 ] = 8'hE8;
  picture_data[ 558 ] = 8'h09;
  picture_data[ 559 ] = 8'hA6;
  picture_data[ 560 ] = 8'h19;
  picture_data[ 561 ] = 8'hC6;
  picture_data[ 562 ] = 8'h09;
  picture_data[ 563 ] = 8'h03;
  picture_data[ 564 ] = 8'h19;
  picture_data[ 565 ] = 8'h04;
  picture_data[ 566 ] = 8'h19;
  picture_data[ 567 ] = 8'h04;
  picture_data[ 568 ] = 8'h21;
  picture_data[ 569 ] = 8'h03;
  picture_data[ 570 ] = 8'h21;
  picture_data[ 571 ] = 8'h02;
  picture_data[ 572 ] = 8'h29;
  picture_data[ 573 ] = 8'h44;
  picture_data[ 574 ] = 8'h29;
  picture_data[ 575 ] = 8'h64;
  picture_data[ 576 ] = 8'h19;
  picture_data[ 577 ] = 8'h83;
  picture_data[ 578 ] = 8'h19;
  picture_data[ 579 ] = 8'h83;
  picture_data[ 580 ] = 8'h29;
  picture_data[ 581 ] = 8'h84;
  picture_data[ 582 ] = 8'h31;
  picture_data[ 583 ] = 8'h84;
  picture_data[ 584 ] = 8'h20;
  picture_data[ 585 ] = 8'hE2;
  picture_data[ 586 ] = 8'h18;
  picture_data[ 587 ] = 8'h80;
  picture_data[ 588 ] = 8'h41;
  picture_data[ 589 ] = 8'hA5;
  picture_data[ 590 ] = 8'h52;
  picture_data[ 591 ] = 8'h47;
  picture_data[ 592 ] = 8'h5A;
  picture_data[ 593 ] = 8'h67;
  picture_data[ 594 ] = 8'h83;
  picture_data[ 595 ] = 8'h8B;
  picture_data[ 596 ] = 8'hBD;
  picture_data[ 597 ] = 8'h52;
  picture_data[ 598 ] = 8'hDE;
  picture_data[ 599 ] = 8'h35;
  picture_data[ 600 ] = 8'hE6;
  picture_data[ 601 ] = 8'h96;
  picture_data[ 602 ] = 8'hD6;
  picture_data[ 603 ] = 8'h13;
  picture_data[ 604 ] = 8'hCD;
  picture_data[ 605 ] = 8'hB1;
  picture_data[ 606 ] = 8'hD6;
  picture_data[ 607 ] = 8'h13;
  picture_data[ 608 ] = 8'h63;
  picture_data[ 609 ] = 8'h2A;
  picture_data[ 610 ] = 8'h21;
  picture_data[ 611 ] = 8'h63;
  picture_data[ 612 ] = 8'h19;
  picture_data[ 613 ] = 8'h02;
  picture_data[ 614 ] = 8'h19;
  picture_data[ 615 ] = 8'h22;
  picture_data[ 616 ] = 8'h11;
  picture_data[ 617 ] = 8'h02;
  picture_data[ 618 ] = 8'h21;
  picture_data[ 619 ] = 8'h63;
  picture_data[ 620 ] = 8'h31;
  picture_data[ 621 ] = 8'hE5;
  picture_data[ 622 ] = 8'h29;
  picture_data[ 623 ] = 8'hA4;
  picture_data[ 624 ] = 8'h5B;
  picture_data[ 625 ] = 8'h09;
  picture_data[ 626 ] = 8'h6B;
  picture_data[ 627 ] = 8'h6B;
  picture_data[ 628 ] = 8'h6B;
  picture_data[ 629 ] = 8'h2A;
  picture_data[ 630 ] = 8'h62;
  picture_data[ 631 ] = 8'hE9;
  picture_data[ 632 ] = 8'h39;
  picture_data[ 633 ] = 8'h84;
  picture_data[ 634 ] = 8'h29;
  picture_data[ 635 ] = 8'h44;
  picture_data[ 636 ] = 8'h31;
  picture_data[ 637 ] = 8'hA6;
  picture_data[ 638 ] = 8'h31;
  picture_data[ 639 ] = 8'hA6;
  picture_data[ 640 ] = 8'h42;
  picture_data[ 641 ] = 8'h47;
  picture_data[ 642 ] = 8'h31;
  picture_data[ 643 ] = 8'hC5;
  picture_data[ 644 ] = 8'h31;
  picture_data[ 645 ] = 8'h43;
  picture_data[ 646 ] = 8'h41;
  picture_data[ 647 ] = 8'hE6;
  picture_data[ 648 ] = 8'h4A;
  picture_data[ 649 ] = 8'h47;
  picture_data[ 650 ] = 8'h63;
  picture_data[ 651 ] = 8'h4B;
  picture_data[ 652 ] = 8'h29;
  picture_data[ 653 ] = 8'hC5;
  picture_data[ 654 ] = 8'h19;
  picture_data[ 655 ] = 8'h64;
  picture_data[ 656 ] = 8'h21;
  picture_data[ 657 ] = 8'h84;
  picture_data[ 658 ] = 8'h19;
  picture_data[ 659 ] = 8'h43;
  picture_data[ 660 ] = 8'h19;
  picture_data[ 661 ] = 8'h23;
  picture_data[ 662 ] = 8'h21;
  picture_data[ 663 ] = 8'h63;
  picture_data[ 664 ] = 8'h29;
  picture_data[ 665 ] = 8'hA4;
  picture_data[ 666 ] = 8'h31;
  picture_data[ 667 ] = 8'hC5;
  picture_data[ 668 ] = 8'h29;
  picture_data[ 669 ] = 8'h64;
  picture_data[ 670 ] = 8'h18;
  picture_data[ 671 ] = 8'hC2;
  picture_data[ 672 ] = 8'h29;
  picture_data[ 673 ] = 8'h64;
  picture_data[ 674 ] = 8'h31;
  picture_data[ 675 ] = 8'h64;
  picture_data[ 676 ] = 8'h20;
  picture_data[ 677 ] = 8'hE2;
  picture_data[ 678 ] = 8'h29;
  picture_data[ 679 ] = 8'h23;
  picture_data[ 680 ] = 8'h31;
  picture_data[ 681 ] = 8'h45;
  picture_data[ 682 ] = 8'h31;
  picture_data[ 683 ] = 8'h04;
  picture_data[ 684 ] = 8'h39;
  picture_data[ 685 ] = 8'h23;
  picture_data[ 686 ] = 8'h28;
  picture_data[ 687 ] = 8'hC1;
  picture_data[ 688 ] = 8'h20;
  picture_data[ 689 ] = 8'hE3;
  picture_data[ 690 ] = 8'h31;
  picture_data[ 691 ] = 8'hC6;
  picture_data[ 692 ] = 8'h29;
  picture_data[ 693 ] = 8'hE7;
  picture_data[ 694 ] = 8'h22;
  picture_data[ 695 ] = 8'h28;
  picture_data[ 696 ] = 8'h1A;
  picture_data[ 697 ] = 8'hAB;
  picture_data[ 698 ] = 8'h23;
  picture_data[ 699 ] = 8'hF0;
  picture_data[ 700 ] = 8'h45;
  picture_data[ 701 ] = 8'hF8;
  picture_data[ 702 ] = 8'h2D;
  picture_data[ 703 ] = 8'h97;
  picture_data[ 704 ] = 8'h03;
  picture_data[ 705 ] = 8'h4D;
  picture_data[ 706 ] = 8'h02;
  picture_data[ 707 ] = 8'h8A;
  picture_data[ 708 ] = 8'h0A;
  picture_data[ 709 ] = 8'h09;
  picture_data[ 710 ] = 8'h01;
  picture_data[ 711 ] = 8'h66;
  picture_data[ 712 ] = 8'h09;
  picture_data[ 713 ] = 8'h44;
  picture_data[ 714 ] = 8'h09;
  picture_data[ 715 ] = 8'h03;
  picture_data[ 716 ] = 8'h10;
  picture_data[ 717 ] = 8'hE3;
  picture_data[ 718 ] = 8'h21;
  picture_data[ 719 ] = 8'h25;
  picture_data[ 720 ] = 8'h10;
  picture_data[ 721 ] = 8'hC3;
  picture_data[ 722 ] = 8'h21;
  picture_data[ 723 ] = 8'h03;
  picture_data[ 724 ] = 8'h29;
  picture_data[ 725 ] = 8'h44;
  picture_data[ 726 ] = 8'h29;
  picture_data[ 727 ] = 8'h64;
  picture_data[ 728 ] = 8'h21;
  picture_data[ 729 ] = 8'h63;
  picture_data[ 730 ] = 8'h21;
  picture_data[ 731 ] = 8'h42;
  picture_data[ 732 ] = 8'h20;
  picture_data[ 733 ] = 8'hE2;
  picture_data[ 734 ] = 8'h31;
  picture_data[ 735 ] = 8'h24;
  picture_data[ 736 ] = 8'h28;
  picture_data[ 737 ] = 8'hE2;
  picture_data[ 738 ] = 8'h39;
  picture_data[ 739 ] = 8'h23;
  picture_data[ 740 ] = 8'h49;
  picture_data[ 741 ] = 8'h84;
  picture_data[ 742 ] = 8'h5A;
  picture_data[ 743 ] = 8'h06;
  picture_data[ 744 ] = 8'h5A;
  picture_data[ 745 ] = 8'h26;
  picture_data[ 746 ] = 8'h7B;
  picture_data[ 747 ] = 8'h09;
  picture_data[ 748 ] = 8'hBD;
  picture_data[ 749 ] = 8'h31;
  picture_data[ 750 ] = 8'hDE;
  picture_data[ 751 ] = 8'h14;
  picture_data[ 752 ] = 8'hDE;
  picture_data[ 753 ] = 8'h13;
  picture_data[ 754 ] = 8'hDE;
  picture_data[ 755 ] = 8'h33;
  picture_data[ 756 ] = 8'hCD;
  picture_data[ 757 ] = 8'hD2;
  picture_data[ 758 ] = 8'hCD;
  picture_data[ 759 ] = 8'hD1;
  picture_data[ 760 ] = 8'h21;
  picture_data[ 761 ] = 8'h42;
  picture_data[ 762 ] = 8'h21;
  picture_data[ 763 ] = 8'h42;
  picture_data[ 764 ] = 8'h21;
  picture_data[ 765 ] = 8'h43;
  picture_data[ 766 ] = 8'h08;
  picture_data[ 767 ] = 8'h80;
  picture_data[ 768 ] = 8'h21;
  picture_data[ 769 ] = 8'h64;
  picture_data[ 770 ] = 8'h29;
  picture_data[ 771 ] = 8'hA5;
  picture_data[ 772 ] = 8'h21;
  picture_data[ 773 ] = 8'h84;
  picture_data[ 774 ] = 8'h29;
  picture_data[ 775 ] = 8'hA4;
  picture_data[ 776 ] = 8'h42;
  picture_data[ 777 ] = 8'h47;
  picture_data[ 778 ] = 8'h39;
  picture_data[ 779 ] = 8'hC5;
  picture_data[ 780 ] = 8'h42;
  picture_data[ 781 ] = 8'h06;
  picture_data[ 782 ] = 8'h41;
  picture_data[ 783 ] = 8'hE6;
  picture_data[ 784 ] = 8'h31;
  picture_data[ 785 ] = 8'h64;
  picture_data[ 786 ] = 8'h31;
  picture_data[ 787 ] = 8'h85;
  picture_data[ 788 ] = 8'h29;
  picture_data[ 789 ] = 8'h65;
  picture_data[ 790 ] = 8'h21;
  picture_data[ 791 ] = 8'h44;
  picture_data[ 792 ] = 8'h29;
  picture_data[ 793 ] = 8'h64;
  picture_data[ 794 ] = 8'h29;
  picture_data[ 795 ] = 8'h64;
  picture_data[ 796 ] = 8'h31;
  picture_data[ 797 ] = 8'h84;
  picture_data[ 798 ] = 8'h39;
  picture_data[ 799 ] = 8'hC5;
  picture_data[ 800 ] = 8'h39;
  picture_data[ 801 ] = 8'hC5;
  picture_data[ 802 ] = 8'h29;
  picture_data[ 803 ] = 8'hA5;
  picture_data[ 804 ] = 8'h19;
  picture_data[ 805 ] = 8'h43;
  picture_data[ 806 ] = 8'h32;
  picture_data[ 807 ] = 8'h06;
  picture_data[ 808 ] = 8'h21;
  picture_data[ 809 ] = 8'h64;
  picture_data[ 810 ] = 8'h19;
  picture_data[ 811 ] = 8'h43;
  picture_data[ 812 ] = 8'h21;
  picture_data[ 813 ] = 8'h43;
  picture_data[ 814 ] = 8'h29;
  picture_data[ 815 ] = 8'h84;
  picture_data[ 816 ] = 8'h21;
  picture_data[ 817 ] = 8'h43;
  picture_data[ 818 ] = 8'h29;
  picture_data[ 819 ] = 8'h64;
  picture_data[ 820 ] = 8'h31;
  picture_data[ 821 ] = 8'h84;
  picture_data[ 822 ] = 8'h31;
  picture_data[ 823 ] = 8'hA5;
  picture_data[ 824 ] = 8'h31;
  picture_data[ 825 ] = 8'h64;
  picture_data[ 826 ] = 8'h31;
  picture_data[ 827 ] = 8'h64;
  picture_data[ 828 ] = 8'h31;
  picture_data[ 829 ] = 8'h23;
  picture_data[ 830 ] = 8'h28;
  picture_data[ 831 ] = 8'hE3;
  picture_data[ 832 ] = 8'h18;
  picture_data[ 833 ] = 8'h21;
  picture_data[ 834 ] = 8'h30;
  picture_data[ 835 ] = 8'hC3;
  picture_data[ 836 ] = 8'h38;
  picture_data[ 837 ] = 8'h81;
  picture_data[ 838 ] = 8'h38;
  picture_data[ 839 ] = 8'hA1;
  picture_data[ 840 ] = 8'h39;
  picture_data[ 841 ] = 8'h23;
  picture_data[ 842 ] = 8'h31;
  picture_data[ 843 ] = 8'h24;
  picture_data[ 844 ] = 8'h29;
  picture_data[ 845 ] = 8'h66;
  picture_data[ 846 ] = 8'h32;
  picture_data[ 847 ] = 8'h29;
  picture_data[ 848 ] = 8'h12;
  picture_data[ 849 ] = 8'h49;
  picture_data[ 850 ] = 8'h0A;
  picture_data[ 851 ] = 8'hAB;
  picture_data[ 852 ] = 8'h02;
  picture_data[ 853 ] = 8'h8B;
  picture_data[ 854 ] = 8'h02;
  picture_data[ 855 ] = 8'h4A;
  picture_data[ 856 ] = 8'h0A;
  picture_data[ 857 ] = 8'hEC;
  picture_data[ 858 ] = 8'h12;
  picture_data[ 859 ] = 8'hAB;
  picture_data[ 860 ] = 8'h1A;
  picture_data[ 861 ] = 8'h4A;
  picture_data[ 862 ] = 8'h11;
  picture_data[ 863 ] = 8'hC8;
  picture_data[ 864 ] = 8'h01;
  picture_data[ 865 ] = 8'h04;
  picture_data[ 866 ] = 8'h11;
  picture_data[ 867 ] = 8'h44;
  picture_data[ 868 ] = 8'h08;
  picture_data[ 869 ] = 8'hC3;
  picture_data[ 870 ] = 8'h19;
  picture_data[ 871 ] = 8'h25;
  picture_data[ 872 ] = 8'h10;
  picture_data[ 873 ] = 8'hC3;
  picture_data[ 874 ] = 8'h19;
  picture_data[ 875 ] = 8'h04;
  picture_data[ 876 ] = 8'h21;
  picture_data[ 877 ] = 8'h24;
  picture_data[ 878 ] = 8'h31;
  picture_data[ 879 ] = 8'h65;
  picture_data[ 880 ] = 8'h18;
  picture_data[ 881 ] = 8'hE2;
  picture_data[ 882 ] = 8'h18;
  picture_data[ 883 ] = 8'hC2;
  picture_data[ 884 ] = 8'h20;
  picture_data[ 885 ] = 8'hC3;
  picture_data[ 886 ] = 8'h39;
  picture_data[ 887 ] = 8'h24;
  picture_data[ 888 ] = 8'h38;
  picture_data[ 889 ] = 8'hE2;
  picture_data[ 890 ] = 8'h6A;
  picture_data[ 891 ] = 8'h27;
  picture_data[ 892 ] = 8'hAC;
  picture_data[ 893 ] = 8'h2F;
  picture_data[ 894 ] = 8'hCD;
  picture_data[ 895 ] = 8'h52;
  picture_data[ 896 ] = 8'hA4;
  picture_data[ 897 ] = 8'h0D;
  picture_data[ 898 ] = 8'h9B;
  picture_data[ 899 ] = 8'hEC;
  picture_data[ 900 ] = 8'hC5;
  picture_data[ 901 ] = 8'h31;
  picture_data[ 902 ] = 8'hC5;
  picture_data[ 903 ] = 8'h51;
  picture_data[ 904 ] = 8'hDE;
  picture_data[ 905 ] = 8'h13;
  picture_data[ 906 ] = 8'hDE;
  picture_data[ 907 ] = 8'h33;
  picture_data[ 908 ] = 8'hDE;
  picture_data[ 909 ] = 8'h13;
  picture_data[ 910 ] = 8'hCD;
  picture_data[ 911 ] = 8'hB1;
  picture_data[ 912 ] = 8'h19;
  picture_data[ 913 ] = 8'h22;
  picture_data[ 914 ] = 8'h3A;
  picture_data[ 915 ] = 8'h06;
  picture_data[ 916 ] = 8'h21;
  picture_data[ 917 ] = 8'h23;
  picture_data[ 918 ] = 8'h21;
  picture_data[ 919 ] = 8'h02;
  picture_data[ 920 ] = 8'h31;
  picture_data[ 921 ] = 8'hA5;
  picture_data[ 922 ] = 8'h21;
  picture_data[ 923 ] = 8'h43;
  picture_data[ 924 ] = 8'h29;
  picture_data[ 925 ] = 8'hC5;
  picture_data[ 926 ] = 8'h3A;
  picture_data[ 927 ] = 8'h47;
  picture_data[ 928 ] = 8'h3A;
  picture_data[ 929 ] = 8'h46;
  picture_data[ 930 ] = 8'h31;
  picture_data[ 931 ] = 8'hE5;
  picture_data[ 932 ] = 8'h39;
  picture_data[ 933 ] = 8'hC5;
  picture_data[ 934 ] = 8'h31;
  picture_data[ 935 ] = 8'h84;
  picture_data[ 936 ] = 8'h39;
  picture_data[ 937 ] = 8'hA5;
  picture_data[ 938 ] = 8'h3A;
  picture_data[ 939 ] = 8'h07;
  picture_data[ 940 ] = 8'h29;
  picture_data[ 941 ] = 8'hA5;
  picture_data[ 942 ] = 8'h21;
  picture_data[ 943 ] = 8'h64;
  picture_data[ 944 ] = 8'h31;
  picture_data[ 945 ] = 8'hC5;
  picture_data[ 946 ] = 8'h29;
  picture_data[ 947 ] = 8'h84;
  picture_data[ 948 ] = 8'h31;
  picture_data[ 949 ] = 8'h84;
  picture_data[ 950 ] = 8'h39;
  picture_data[ 951 ] = 8'hA5;
  picture_data[ 952 ] = 8'h39;
  picture_data[ 953 ] = 8'hC5;
  picture_data[ 954 ] = 8'h19;
  picture_data[ 955 ] = 8'h02;
  picture_data[ 956 ] = 8'h21;
  picture_data[ 957 ] = 8'h63;
  picture_data[ 958 ] = 8'h29;
  picture_data[ 959 ] = 8'h85;
  picture_data[ 960 ] = 8'h19;
  picture_data[ 961 ] = 8'h43;
  picture_data[ 962 ] = 8'h19;
  picture_data[ 963 ] = 8'h02;
  picture_data[ 964 ] = 8'h10;
  picture_data[ 965 ] = 8'hE2;
  picture_data[ 966 ] = 8'h31;
  picture_data[ 967 ] = 8'hC5;
  picture_data[ 968 ] = 8'h39;
  picture_data[ 969 ] = 8'hC5;
  picture_data[ 970 ] = 8'h31;
  picture_data[ 971 ] = 8'h84;
  picture_data[ 972 ] = 8'h31;
  picture_data[ 973 ] = 8'h64;
  picture_data[ 974 ] = 8'h4A;
  picture_data[ 975 ] = 8'h47;
  picture_data[ 976 ] = 8'h21;
  picture_data[ 977 ] = 8'h02;
  picture_data[ 978 ] = 8'h29;
  picture_data[ 979 ] = 8'h23;
  picture_data[ 980 ] = 8'h39;
  picture_data[ 981 ] = 8'h44;
  picture_data[ 982 ] = 8'h30;
  picture_data[ 983 ] = 8'hC3;
  picture_data[ 984 ] = 8'h28;
  picture_data[ 985 ] = 8'h63;
  picture_data[ 986 ] = 8'h30;
  picture_data[ 987 ] = 8'h22;
  picture_data[ 988 ] = 8'h50;
  picture_data[ 989 ] = 8'h82;
  picture_data[ 990 ] = 8'h58;
  picture_data[ 991 ] = 8'hA2;
  picture_data[ 992 ] = 8'h58;
  picture_data[ 993 ] = 8'hA2;
  picture_data[ 994 ] = 8'h59;
  picture_data[ 995 ] = 8'h04;
  picture_data[ 996 ] = 8'h51;
  picture_data[ 997 ] = 8'h05;
  picture_data[ 998 ] = 8'h41;
  picture_data[ 999 ] = 8'h67;
  picture_data[ 1000 ] = 8'h19;
  picture_data[ 1001 ] = 8'hC8;
  picture_data[ 1002 ] = 8'h22;
  picture_data[ 1003 ] = 8'hCC;
  picture_data[ 1004 ] = 8'h22;
  picture_data[ 1005 ] = 8'h6A;
  picture_data[ 1006 ] = 8'h09;
  picture_data[ 1007 ] = 8'hC7;
  picture_data[ 1008 ] = 8'h23;
  picture_data[ 1009 ] = 8'h0D;
  picture_data[ 1010 ] = 8'h22;
  picture_data[ 1011 ] = 8'hCC;
  picture_data[ 1012 ] = 8'h01;
  picture_data[ 1013 ] = 8'h46;
  picture_data[ 1014 ] = 8'h11;
  picture_data[ 1015 ] = 8'h87;
  picture_data[ 1016 ] = 8'h09;
  picture_data[ 1017 ] = 8'h46;
  picture_data[ 1018 ] = 8'h01;
  picture_data[ 1019 ] = 8'h04;
  picture_data[ 1020 ] = 8'h19;
  picture_data[ 1021 ] = 8'h87;
  picture_data[ 1022 ] = 8'h19;
  picture_data[ 1023 ] = 8'h66;
  picture_data[ 1024 ] = 8'h19;
  picture_data[ 1025 ] = 8'h45;
  picture_data[ 1026 ] = 8'h19;
  picture_data[ 1027 ] = 8'h04;
  picture_data[ 1028 ] = 8'h21;
  picture_data[ 1029 ] = 8'h24;
  picture_data[ 1030 ] = 8'h31;
  picture_data[ 1031 ] = 8'h85;
  picture_data[ 1032 ] = 8'h31;
  picture_data[ 1033 ] = 8'hA6;
  picture_data[ 1034 ] = 8'h29;
  picture_data[ 1035 ] = 8'h44;
  picture_data[ 1036 ] = 8'h39;
  picture_data[ 1037 ] = 8'h65;
  picture_data[ 1038 ] = 8'h41;
  picture_data[ 1039 ] = 8'h04;
  picture_data[ 1040 ] = 8'h59;
  picture_data[ 1041 ] = 8'h43;
  picture_data[ 1042 ] = 8'h8A;
  picture_data[ 1043 ] = 8'hC9;
  picture_data[ 1044 ] = 8'hAB;
  picture_data[ 1045 ] = 8'hCC;
  picture_data[ 1046 ] = 8'hDD;
  picture_data[ 1047 ] = 8'h73;
  picture_data[ 1048 ] = 8'hFE;
  picture_data[ 1049 ] = 8'hB7;
  picture_data[ 1050 ] = 8'hEE;
  picture_data[ 1051 ] = 8'h55;
  picture_data[ 1052 ] = 8'hEE;
  picture_data[ 1053 ] = 8'h75;
  picture_data[ 1054 ] = 8'hE6;
  picture_data[ 1055 ] = 8'h75;
  picture_data[ 1056 ] = 8'hE6;
  picture_data[ 1057 ] = 8'h54;
  picture_data[ 1058 ] = 8'hD5;
  picture_data[ 1059 ] = 8'hF2;
  picture_data[ 1060 ] = 8'hDE;
  picture_data[ 1061 ] = 8'h33;
  picture_data[ 1062 ] = 8'hD6;
  picture_data[ 1063 ] = 8'h12;
  picture_data[ 1064 ] = 8'h3A;
  picture_data[ 1065 ] = 8'h06;
  picture_data[ 1066 ] = 8'h42;
  picture_data[ 1067 ] = 8'h26;
  picture_data[ 1068 ] = 8'h21;
  picture_data[ 1069 ] = 8'h22;
  picture_data[ 1070 ] = 8'h42;
  picture_data[ 1071 ] = 8'h06;
  picture_data[ 1072 ] = 8'h39;
  picture_data[ 1073 ] = 8'hC5;
  picture_data[ 1074 ] = 8'h21;
  picture_data[ 1075 ] = 8'h43;
  picture_data[ 1076 ] = 8'h29;
  picture_data[ 1077 ] = 8'hA5;
  picture_data[ 1078 ] = 8'h52;
  picture_data[ 1079 ] = 8'hE9;
  picture_data[ 1080 ] = 8'h42;
  picture_data[ 1081 ] = 8'h67;
  picture_data[ 1082 ] = 8'h29;
  picture_data[ 1083 ] = 8'h84;
  picture_data[ 1084 ] = 8'h21;
  picture_data[ 1085 ] = 8'h22;
  picture_data[ 1086 ] = 8'h31;
  picture_data[ 1087 ] = 8'h84;
  picture_data[ 1088 ] = 8'h29;
  picture_data[ 1089 ] = 8'h84;
  picture_data[ 1090 ] = 8'h21;
  picture_data[ 1091 ] = 8'h23;
  picture_data[ 1092 ] = 8'h19;
  picture_data[ 1093 ] = 8'h43;
  picture_data[ 1094 ] = 8'h21;
  picture_data[ 1095 ] = 8'h84;
  picture_data[ 1096 ] = 8'h29;
  picture_data[ 1097 ] = 8'hA4;
  picture_data[ 1098 ] = 8'h31;
  picture_data[ 1099 ] = 8'h84;
  picture_data[ 1100 ] = 8'h21;
  picture_data[ 1101 ] = 8'h23;
  picture_data[ 1102 ] = 8'h39;
  picture_data[ 1103 ] = 8'hE5;
  picture_data[ 1104 ] = 8'h21;
  picture_data[ 1105 ] = 8'h23;
  picture_data[ 1106 ] = 8'h21;
  picture_data[ 1107 ] = 8'h23;
  picture_data[ 1108 ] = 8'h19;
  picture_data[ 1109 ] = 8'h02;
  picture_data[ 1110 ] = 8'h10;
  picture_data[ 1111 ] = 8'hE2;
  picture_data[ 1112 ] = 8'h11;
  picture_data[ 1113 ] = 8'h02;
  picture_data[ 1114 ] = 8'h21;
  picture_data[ 1115 ] = 8'h64;
  picture_data[ 1116 ] = 8'h29;
  picture_data[ 1117 ] = 8'h84;
  picture_data[ 1118 ] = 8'h21;
  picture_data[ 1119 ] = 8'h43;
  picture_data[ 1120 ] = 8'h39;
  picture_data[ 1121 ] = 8'hC5;
  picture_data[ 1122 ] = 8'h63;
  picture_data[ 1123 ] = 8'h0A;
  picture_data[ 1124 ] = 8'h4A;
  picture_data[ 1125 ] = 8'h26;
  picture_data[ 1126 ] = 8'h31;
  picture_data[ 1127 ] = 8'h84;
  picture_data[ 1128 ] = 8'h31;
  picture_data[ 1129 ] = 8'h64;
  picture_data[ 1130 ] = 8'h21;
  picture_data[ 1131 ] = 8'h02;
  picture_data[ 1132 ] = 8'h20;
  picture_data[ 1133 ] = 8'h81;
  picture_data[ 1134 ] = 8'h28;
  picture_data[ 1135 ] = 8'h61;
  picture_data[ 1136 ] = 8'h30;
  picture_data[ 1137 ] = 8'h42;
  picture_data[ 1138 ] = 8'h48;
  picture_data[ 1139 ] = 8'hA4;
  picture_data[ 1140 ] = 8'h71;
  picture_data[ 1141 ] = 8'h05;
  picture_data[ 1142 ] = 8'hA2;
  picture_data[ 1143 ] = 8'h4A;
  picture_data[ 1144 ] = 8'hD3;
  picture_data[ 1145 ] = 8'hEF;
  picture_data[ 1146 ] = 8'hC3;
  picture_data[ 1147 ] = 8'h8E;
  picture_data[ 1148 ] = 8'h81;
  picture_data[ 1149 ] = 8'h88;
  picture_data[ 1150 ] = 8'h50;
  picture_data[ 1151 ] = 8'hE6;
  picture_data[ 1152 ] = 8'h29;
  picture_data[ 1153 ] = 8'hA9;
  picture_data[ 1154 ] = 8'h22;
  picture_data[ 1155 ] = 8'h0B;
  picture_data[ 1156 ] = 8'h29;
  picture_data[ 1157 ] = 8'hE9;
  picture_data[ 1158 ] = 8'h21;
  picture_data[ 1159 ] = 8'hA8;
  picture_data[ 1160 ] = 8'h12;
  picture_data[ 1161 ] = 8'h0A;
  picture_data[ 1162 ] = 8'h12;
  picture_data[ 1163 ] = 8'h2A;
  picture_data[ 1164 ] = 8'h11;
  picture_data[ 1165 ] = 8'hA9;
  picture_data[ 1166 ] = 8'h09;
  picture_data[ 1167 ] = 8'h26;
  picture_data[ 1168 ] = 8'h09;
  picture_data[ 1169 ] = 8'h26;
  picture_data[ 1170 ] = 8'h11;
  picture_data[ 1171 ] = 8'h26;
  picture_data[ 1172 ] = 8'h11;
  picture_data[ 1173 ] = 8'h05;
  picture_data[ 1174 ] = 8'h21;
  picture_data[ 1175 ] = 8'h66;
  picture_data[ 1176 ] = 8'h21;
  picture_data[ 1177 ] = 8'h45;
  picture_data[ 1178 ] = 8'h21;
  picture_data[ 1179 ] = 8'h25;
  picture_data[ 1180 ] = 8'h29;
  picture_data[ 1181 ] = 8'h65;
  picture_data[ 1182 ] = 8'h31;
  picture_data[ 1183 ] = 8'h85;
  picture_data[ 1184 ] = 8'h73;
  picture_data[ 1185 ] = 8'h8D;
  picture_data[ 1186 ] = 8'h5A;
  picture_data[ 1187 ] = 8'hA9;
  picture_data[ 1188 ] = 8'h73;
  picture_data[ 1189 ] = 8'h2B;
  picture_data[ 1190 ] = 8'h83;
  picture_data[ 1191 ] = 8'h2B;
  picture_data[ 1192 ] = 8'h72;
  picture_data[ 1193 ] = 8'h26;
  picture_data[ 1194 ] = 8'hFE;
  picture_data[ 1195 ] = 8'h77;
  picture_data[ 1196 ] = 8'hED;
  picture_data[ 1197 ] = 8'hD4;
  picture_data[ 1198 ] = 8'hBC;
  picture_data[ 1199 ] = 8'h8F;
  picture_data[ 1200 ] = 8'hF6;
  picture_data[ 1201 ] = 8'h56;
  picture_data[ 1202 ] = 8'hEE;
  picture_data[ 1203 ] = 8'h55;
  picture_data[ 1204 ] = 8'hE6;
  picture_data[ 1205 ] = 8'h34;
  picture_data[ 1206 ] = 8'hDE;
  picture_data[ 1207 ] = 8'h54;
  picture_data[ 1208 ] = 8'hDE;
  picture_data[ 1209 ] = 8'h34;
  picture_data[ 1210 ] = 8'hDE;
  picture_data[ 1211 ] = 8'h54;
  picture_data[ 1212 ] = 8'hDE;
  picture_data[ 1213 ] = 8'h33;
  picture_data[ 1214 ] = 8'hD6;
  picture_data[ 1215 ] = 8'h13;
  picture_data[ 1216 ] = 8'h21;
  picture_data[ 1217 ] = 8'h02;
  picture_data[ 1218 ] = 8'h29;
  picture_data[ 1219 ] = 8'h63;
  picture_data[ 1220 ] = 8'h31;
  picture_data[ 1221 ] = 8'h84;
  picture_data[ 1222 ] = 8'h83;
  picture_data[ 1223 ] = 8'hED;
  picture_data[ 1224 ] = 8'h39;
  picture_data[ 1225 ] = 8'hA5;
  picture_data[ 1226 ] = 8'h21;
  picture_data[ 1227 ] = 8'h43;
  picture_data[ 1228 ] = 8'h21;
  picture_data[ 1229 ] = 8'h63;
  picture_data[ 1230 ] = 8'h19;
  picture_data[ 1231 ] = 8'h43;
  picture_data[ 1232 ] = 8'h21;
  picture_data[ 1233 ] = 8'h63;
  picture_data[ 1234 ] = 8'h3A;
  picture_data[ 1235 ] = 8'h06;
  picture_data[ 1236 ] = 8'h42;
  picture_data[ 1237 ] = 8'h46;
  picture_data[ 1238 ] = 8'h31;
  picture_data[ 1239 ] = 8'hA4;
  picture_data[ 1240 ] = 8'h29;
  picture_data[ 1241 ] = 8'h84;
  picture_data[ 1242 ] = 8'h29;
  picture_data[ 1243 ] = 8'hA4;
  picture_data[ 1244 ] = 8'h21;
  picture_data[ 1245 ] = 8'h63;
  picture_data[ 1246 ] = 8'h19;
  picture_data[ 1247 ] = 8'h63;
  picture_data[ 1248 ] = 8'h29;
  picture_data[ 1249 ] = 8'hA4;
  picture_data[ 1250 ] = 8'h29;
  picture_data[ 1251 ] = 8'h63;
  picture_data[ 1252 ] = 8'h21;
  picture_data[ 1253 ] = 8'h43;
  picture_data[ 1254 ] = 8'h21;
  picture_data[ 1255 ] = 8'h23;
  picture_data[ 1256 ] = 8'h18;
  picture_data[ 1257 ] = 8'hE2;
  picture_data[ 1258 ] = 8'h19;
  picture_data[ 1259 ] = 8'h02;
  picture_data[ 1260 ] = 8'h19;
  picture_data[ 1261 ] = 8'h23;
  picture_data[ 1262 ] = 8'h21;
  picture_data[ 1263 ] = 8'h44;
  picture_data[ 1264 ] = 8'h19;
  picture_data[ 1265 ] = 8'h23;
  picture_data[ 1266 ] = 8'h19;
  picture_data[ 1267 ] = 8'h43;
  picture_data[ 1268 ] = 8'h21;
  picture_data[ 1269 ] = 8'h84;
  picture_data[ 1270 ] = 8'h29;
  picture_data[ 1271 ] = 8'hA5;
  picture_data[ 1272 ] = 8'h29;
  picture_data[ 1273 ] = 8'h63;
  picture_data[ 1274 ] = 8'h4A;
  picture_data[ 1275 ] = 8'h88;
  picture_data[ 1276 ] = 8'h4A;
  picture_data[ 1277 ] = 8'h67;
  picture_data[ 1278 ] = 8'h21;
  picture_data[ 1279 ] = 8'h02;
  picture_data[ 1280 ] = 8'h29;
  picture_data[ 1281 ] = 8'h23;
  picture_data[ 1282 ] = 8'h20;
  picture_data[ 1283 ] = 8'hE2;
  picture_data[ 1284 ] = 8'h20;
  picture_data[ 1285 ] = 8'hA0;
  picture_data[ 1286 ] = 8'h39;
  picture_data[ 1287 ] = 8'h23;
  picture_data[ 1288 ] = 8'h51;
  picture_data[ 1289 ] = 8'h85;
  picture_data[ 1290 ] = 8'h71;
  picture_data[ 1291 ] = 8'hE7;
  picture_data[ 1292 ] = 8'h99;
  picture_data[ 1293 ] = 8'hE9;
  picture_data[ 1294 ] = 8'hFE;
  picture_data[ 1295 ] = 8'h5A;
  picture_data[ 1296 ] = 8'hFF;
  picture_data[ 1297 ] = 8'h3C;
  picture_data[ 1298 ] = 8'hFE;
  picture_data[ 1299 ] = 8'h99;
  picture_data[ 1300 ] = 8'hE4;
  picture_data[ 1301 ] = 8'h72;
  picture_data[ 1302 ] = 8'h58;
  picture_data[ 1303 ] = 8'h85;
  picture_data[ 1304 ] = 8'h41;
  picture_data[ 1305 ] = 8'h4B;
  picture_data[ 1306 ] = 8'h21;
  picture_data[ 1307 ] = 8'h4C;
  picture_data[ 1308 ] = 8'h21;
  picture_data[ 1309 ] = 8'h0A;
  picture_data[ 1310 ] = 8'h31;
  picture_data[ 1311 ] = 8'hCC;
  picture_data[ 1312 ] = 8'h22;
  picture_data[ 1313 ] = 8'h2C;
  picture_data[ 1314 ] = 8'h09;
  picture_data[ 1315 ] = 8'hA9;
  picture_data[ 1316 ] = 8'h01;
  picture_data[ 1317 ] = 8'h48;
  picture_data[ 1318 ] = 8'h09;
  picture_data[ 1319 ] = 8'h47;
  picture_data[ 1320 ] = 8'h19;
  picture_data[ 1321 ] = 8'h48;
  picture_data[ 1322 ] = 8'h10;
  picture_data[ 1323 ] = 8'hC5;
  picture_data[ 1324 ] = 8'h18;
  picture_data[ 1325 ] = 8'hC4;
  picture_data[ 1326 ] = 8'h31;
  picture_data[ 1327 ] = 8'h25;
  picture_data[ 1328 ] = 8'h31;
  picture_data[ 1329 ] = 8'h65;
  picture_data[ 1330 ] = 8'h29;
  picture_data[ 1331 ] = 8'h23;
  picture_data[ 1332 ] = 8'h39;
  picture_data[ 1333 ] = 8'hC5;
  picture_data[ 1334 ] = 8'h29;
  picture_data[ 1335 ] = 8'h22;
  picture_data[ 1336 ] = 8'h4A;
  picture_data[ 1337 ] = 8'h06;
  picture_data[ 1338 ] = 8'h83;
  picture_data[ 1339 ] = 8'hED;
  picture_data[ 1340 ] = 8'hBD;
  picture_data[ 1341 ] = 8'hD4;
  picture_data[ 1342 ] = 8'hDE;
  picture_data[ 1343 ] = 8'h77;
  picture_data[ 1344 ] = 8'hF6;
  picture_data[ 1345 ] = 8'h77;
  picture_data[ 1346 ] = 8'hDD;
  picture_data[ 1347 ] = 8'h52;
  picture_data[ 1348 ] = 8'hE5;
  picture_data[ 1349 ] = 8'h93;
  picture_data[ 1350 ] = 8'hE5;
  picture_data[ 1351 ] = 8'hF4;
  picture_data[ 1352 ] = 8'hEE;
  picture_data[ 1353 ] = 8'h55;
  picture_data[ 1354 ] = 8'hE6;
  picture_data[ 1355 ] = 8'h55;
  picture_data[ 1356 ] = 8'hE6;
  picture_data[ 1357 ] = 8'h75;
  picture_data[ 1358 ] = 8'hDE;
  picture_data[ 1359 ] = 8'h54;
  picture_data[ 1360 ] = 8'hDE;
  picture_data[ 1361 ] = 8'h54;
  picture_data[ 1362 ] = 8'hDE;
  picture_data[ 1363 ] = 8'h54;
  picture_data[ 1364 ] = 8'hD6;
  picture_data[ 1365 ] = 8'h33;
  picture_data[ 1366 ] = 8'hD6;
  picture_data[ 1367 ] = 8'h34;
  picture_data[ 1368 ] = 8'h20;
  picture_data[ 1369 ] = 8'hE1;
  picture_data[ 1370 ] = 8'h31;
  picture_data[ 1371 ] = 8'h83;
  picture_data[ 1372 ] = 8'h29;
  picture_data[ 1373 ] = 8'h02;
  picture_data[ 1374 ] = 8'h10;
  picture_data[ 1375 ] = 8'h40;
  picture_data[ 1376 ] = 8'h21;
  picture_data[ 1377 ] = 8'h02;
  picture_data[ 1378 ] = 8'h29;
  picture_data[ 1379 ] = 8'h43;
  picture_data[ 1380 ] = 8'h19;
  picture_data[ 1381 ] = 8'h22;
  picture_data[ 1382 ] = 8'h21;
  picture_data[ 1383 ] = 8'h63;
  picture_data[ 1384 ] = 8'h29;
  picture_data[ 1385 ] = 8'hA4;
  picture_data[ 1386 ] = 8'h19;
  picture_data[ 1387 ] = 8'h42;
  picture_data[ 1388 ] = 8'h29;
  picture_data[ 1389 ] = 8'h63;
  picture_data[ 1390 ] = 8'h21;
  picture_data[ 1391 ] = 8'h22;
  picture_data[ 1392 ] = 8'h19;
  picture_data[ 1393 ] = 8'h02;
  picture_data[ 1394 ] = 8'h31;
  picture_data[ 1395 ] = 8'hC5;
  picture_data[ 1396 ] = 8'h3A;
  picture_data[ 1397 ] = 8'h47;
  picture_data[ 1398 ] = 8'h21;
  picture_data[ 1399 ] = 8'h84;
  picture_data[ 1400 ] = 8'h29;
  picture_data[ 1401 ] = 8'h84;
  picture_data[ 1402 ] = 8'h29;
  picture_data[ 1403 ] = 8'hA4;
  picture_data[ 1404 ] = 8'h32;
  picture_data[ 1405 ] = 8'h06;
  picture_data[ 1406 ] = 8'h29;
  picture_data[ 1407 ] = 8'hC6;
  picture_data[ 1408 ] = 8'h19;
  picture_data[ 1409 ] = 8'h44;
  picture_data[ 1410 ] = 8'h19;
  picture_data[ 1411 ] = 8'h23;
  picture_data[ 1412 ] = 8'h21;
  picture_data[ 1413 ] = 8'h64;
  picture_data[ 1414 ] = 8'h19;
  picture_data[ 1415 ] = 8'h43;
  picture_data[ 1416 ] = 8'h21;
  picture_data[ 1417 ] = 8'hA5;
  picture_data[ 1418 ] = 8'h11;
  picture_data[ 1419 ] = 8'h23;
  picture_data[ 1420 ] = 8'h11;
  picture_data[ 1421 ] = 8'h23;
  picture_data[ 1422 ] = 8'h29;
  picture_data[ 1423 ] = 8'hA5;
  picture_data[ 1424 ] = 8'h19;
  picture_data[ 1425 ] = 8'h43;
  picture_data[ 1426 ] = 8'h21;
  picture_data[ 1427 ] = 8'h64;
  picture_data[ 1428 ] = 8'h21;
  picture_data[ 1429 ] = 8'h43;
  picture_data[ 1430 ] = 8'h21;
  picture_data[ 1431 ] = 8'h02;
  picture_data[ 1432 ] = 8'h18;
  picture_data[ 1433 ] = 8'hE2;
  picture_data[ 1434 ] = 8'h29;
  picture_data[ 1435 ] = 8'h23;
  picture_data[ 1436 ] = 8'h29;
  picture_data[ 1437 ] = 8'h22;
  picture_data[ 1438 ] = 8'h31;
  picture_data[ 1439 ] = 8'h22;
  picture_data[ 1440 ] = 8'h51;
  picture_data[ 1441 ] = 8'hC5;
  picture_data[ 1442 ] = 8'h69;
  picture_data[ 1443 ] = 8'hE7;
  picture_data[ 1444 ] = 8'h9A;
  picture_data[ 1445 ] = 8'h2A;
  picture_data[ 1446 ] = 8'hFD;
  picture_data[ 1447 ] = 8'h36;
  picture_data[ 1448 ] = 8'hFD;
  picture_data[ 1449 ] = 8'h34;
  picture_data[ 1450 ] = 8'hE4;
  picture_data[ 1451 ] = 8'hB2;
  picture_data[ 1452 ] = 8'hCB;
  picture_data[ 1453 ] = 8'h8F;
  picture_data[ 1454 ] = 8'h71;
  picture_data[ 1455 ] = 8'hAA;
  picture_data[ 1456 ] = 8'h39;
  picture_data[ 1457 ] = 8'h6E;
  picture_data[ 1458 ] = 8'h08;
  picture_data[ 1459 ] = 8'hCD;
  picture_data[ 1460 ] = 8'h11;
  picture_data[ 1461 ] = 8'h4F;
  picture_data[ 1462 ] = 8'h11;
  picture_data[ 1463 ] = 8'h6D;
  picture_data[ 1464 ] = 8'h11;
  picture_data[ 1465 ] = 8'hAC;
  picture_data[ 1466 ] = 8'h09;
  picture_data[ 1467 ] = 8'h29;
  picture_data[ 1468 ] = 8'h09;
  picture_data[ 1469 ] = 8'h48;
  picture_data[ 1470 ] = 8'h11;
  picture_data[ 1471 ] = 8'h48;
  picture_data[ 1472 ] = 8'h21;
  picture_data[ 1473 ] = 8'h46;
  picture_data[ 1474 ] = 8'h4A;
  picture_data[ 1475 ] = 8'h29;
  picture_data[ 1476 ] = 8'h5A;
  picture_data[ 1477 ] = 8'h4A;
  picture_data[ 1478 ] = 8'h41;
  picture_data[ 1479 ] = 8'hA5;
  picture_data[ 1480 ] = 8'h49;
  picture_data[ 1481 ] = 8'hA3;
  picture_data[ 1482 ] = 8'h41;
  picture_data[ 1483 ] = 8'hA2;
  picture_data[ 1484 ] = 8'h62;
  picture_data[ 1485 ] = 8'h87;
  picture_data[ 1486 ] = 8'hBD;
  picture_data[ 1487 ] = 8'h93;
  picture_data[ 1488 ] = 8'hE6;
  picture_data[ 1489 ] = 8'hF9;
  picture_data[ 1490 ] = 8'hB5;
  picture_data[ 1491 ] = 8'h72;
  picture_data[ 1492 ] = 8'hBD;
  picture_data[ 1493 ] = 8'hB3;
  picture_data[ 1494 ] = 8'hF7;
  picture_data[ 1495 ] = 8'h5A;
  picture_data[ 1496 ] = 8'hFF;
  picture_data[ 1497 ] = 8'h3A;
  picture_data[ 1498 ] = 8'hEE;
  picture_data[ 1499 ] = 8'h56;
  picture_data[ 1500 ] = 8'hE5;
  picture_data[ 1501 ] = 8'hF4;
  picture_data[ 1502 ] = 8'hEE;
  picture_data[ 1503 ] = 8'h76;
  picture_data[ 1504 ] = 8'hE6;
  picture_data[ 1505 ] = 8'h55;
  picture_data[ 1506 ] = 8'hEE;
  picture_data[ 1507 ] = 8'hB6;
  picture_data[ 1508 ] = 8'hE6;
  picture_data[ 1509 ] = 8'h75;
  picture_data[ 1510 ] = 8'hDE;
  picture_data[ 1511 ] = 8'h75;
  picture_data[ 1512 ] = 8'hDE;
  picture_data[ 1513 ] = 8'h74;
  picture_data[ 1514 ] = 8'hDE;
  picture_data[ 1515 ] = 8'h74;
  picture_data[ 1516 ] = 8'hD6;
  picture_data[ 1517 ] = 8'h54;
  picture_data[ 1518 ] = 8'hD6;
  picture_data[ 1519 ] = 8'h33;
  picture_data[ 1520 ] = 8'h10;
  picture_data[ 1521 ] = 8'h60;
  picture_data[ 1522 ] = 8'h63;
  picture_data[ 1523 ] = 8'h09;
  picture_data[ 1524 ] = 8'h9C;
  picture_data[ 1525 ] = 8'hB0;
  picture_data[ 1526 ] = 8'h18;
  picture_data[ 1527 ] = 8'hA0;
  picture_data[ 1528 ] = 8'h39;
  picture_data[ 1529 ] = 8'hA4;
  picture_data[ 1530 ] = 8'h21;
  picture_data[ 1531 ] = 8'h01;
  picture_data[ 1532 ] = 8'h21;
  picture_data[ 1533 ] = 8'h22;
  picture_data[ 1534 ] = 8'h19;
  picture_data[ 1535 ] = 8'h22;
  picture_data[ 1536 ] = 8'h19;
  picture_data[ 1537 ] = 8'h01;
  picture_data[ 1538 ] = 8'h10;
  picture_data[ 1539 ] = 8'hE1;
  picture_data[ 1540 ] = 8'h10;
  picture_data[ 1541 ] = 8'hE1;
  picture_data[ 1542 ] = 8'h10;
  picture_data[ 1543 ] = 8'hE1;
  picture_data[ 1544 ] = 8'h19;
  picture_data[ 1545 ] = 8'h02;
  picture_data[ 1546 ] = 8'h18;
  picture_data[ 1547 ] = 8'hE2;
  picture_data[ 1548 ] = 8'h21;
  picture_data[ 1549 ] = 8'h63;
  picture_data[ 1550 ] = 8'h29;
  picture_data[ 1551 ] = 8'hA4;
  picture_data[ 1552 ] = 8'h21;
  picture_data[ 1553 ] = 8'h84;
  picture_data[ 1554 ] = 8'h21;
  picture_data[ 1555 ] = 8'h85;
  picture_data[ 1556 ] = 8'h19;
  picture_data[ 1557 ] = 8'h64;
  picture_data[ 1558 ] = 8'h11;
  picture_data[ 1559 ] = 8'h44;
  picture_data[ 1560 ] = 8'h21;
  picture_data[ 1561 ] = 8'hC6;
  picture_data[ 1562 ] = 8'h29;
  picture_data[ 1563 ] = 8'hC6;
  picture_data[ 1564 ] = 8'h29;
  picture_data[ 1565 ] = 8'hC6;
  picture_data[ 1566 ] = 8'h21;
  picture_data[ 1567 ] = 8'hA5;
  picture_data[ 1568 ] = 8'h19;
  picture_data[ 1569 ] = 8'h65;
  picture_data[ 1570 ] = 8'h21;
  picture_data[ 1571 ] = 8'hC6;
  picture_data[ 1572 ] = 8'h19;
  picture_data[ 1573 ] = 8'h85;
  picture_data[ 1574 ] = 8'h19;
  picture_data[ 1575 ] = 8'h65;
  picture_data[ 1576 ] = 8'h11;
  picture_data[ 1577 ] = 8'h03;
  picture_data[ 1578 ] = 8'h19;
  picture_data[ 1579 ] = 8'h23;
  picture_data[ 1580 ] = 8'h11;
  picture_data[ 1581 ] = 8'h03;
  picture_data[ 1582 ] = 8'h19;
  picture_data[ 1583 ] = 8'h02;
  picture_data[ 1584 ] = 8'h19;
  picture_data[ 1585 ] = 8'h03;
  picture_data[ 1586 ] = 8'h29;
  picture_data[ 1587 ] = 8'h44;
  picture_data[ 1588 ] = 8'h31;
  picture_data[ 1589 ] = 8'h44;
  picture_data[ 1590 ] = 8'h30;
  picture_data[ 1591 ] = 8'hE2;
  picture_data[ 1592 ] = 8'h30;
  picture_data[ 1593 ] = 8'hC2;
  picture_data[ 1594 ] = 8'h59;
  picture_data[ 1595 ] = 8'h65;
  picture_data[ 1596 ] = 8'h81;
  picture_data[ 1597 ] = 8'hA8;
  picture_data[ 1598 ] = 8'h89;
  picture_data[ 1599 ] = 8'h88;
  picture_data[ 1600 ] = 8'hA2;
  picture_data[ 1601 ] = 8'h09;
  picture_data[ 1602 ] = 8'h99;
  picture_data[ 1603 ] = 8'hC8;
  picture_data[ 1604 ] = 8'h79;
  picture_data[ 1605 ] = 8'hC8;
  picture_data[ 1606 ] = 8'h59;
  picture_data[ 1607 ] = 8'hEC;
  picture_data[ 1608 ] = 8'h11;
  picture_data[ 1609 ] = 8'h30;
  picture_data[ 1610 ] = 8'h2A;
  picture_data[ 1611 ] = 8'hF9;
  picture_data[ 1612 ] = 8'h34;
  picture_data[ 1613 ] = 8'h1D;
  picture_data[ 1614 ] = 8'h1B;
  picture_data[ 1615 ] = 8'h58;
  picture_data[ 1616 ] = 8'h09;
  picture_data[ 1617 ] = 8'hAF;
  picture_data[ 1618 ] = 8'h09;
  picture_data[ 1619 ] = 8'h0A;
  picture_data[ 1620 ] = 8'h21;
  picture_data[ 1621 ] = 8'h69;
  picture_data[ 1622 ] = 8'h5B;
  picture_data[ 1623 ] = 8'h0D;
  picture_data[ 1624 ] = 8'h5A;
  picture_data[ 1625 ] = 8'hCA;
  picture_data[ 1626 ] = 8'h83;
  picture_data[ 1627 ] = 8'hCE;
  picture_data[ 1628 ] = 8'h62;
  picture_data[ 1629 ] = 8'hC9;
  picture_data[ 1630 ] = 8'h7B;
  picture_data[ 1631 ] = 8'h29;
  picture_data[ 1632 ] = 8'hC5;
  picture_data[ 1633 ] = 8'h0B;
  picture_data[ 1634 ] = 8'hD5;
  picture_data[ 1635 ] = 8'hAD;
  picture_data[ 1636 ] = 8'hE6;
  picture_data[ 1637 ] = 8'h73;
  picture_data[ 1638 ] = 8'hFF;
  picture_data[ 1639 ] = 8'hDC;
  picture_data[ 1640 ] = 8'hFF;
  picture_data[ 1641 ] = 8'hFE;
  picture_data[ 1642 ] = 8'hF7;
  picture_data[ 1643 ] = 8'h9D;
  picture_data[ 1644 ] = 8'hF7;
  picture_data[ 1645 ] = 8'h7C;
  picture_data[ 1646 ] = 8'hF7;
  picture_data[ 1647 ] = 8'h3B;
  picture_data[ 1648 ] = 8'hFF;
  picture_data[ 1649 ] = 8'h7B;
  picture_data[ 1650 ] = 8'hF7;
  picture_data[ 1651 ] = 8'h39;
  picture_data[ 1652 ] = 8'hF7;
  picture_data[ 1653 ] = 8'h19;
  picture_data[ 1654 ] = 8'hEE;
  picture_data[ 1655 ] = 8'hD8;
  picture_data[ 1656 ] = 8'hEE;
  picture_data[ 1657 ] = 8'hD7;
  picture_data[ 1658 ] = 8'hE6;
  picture_data[ 1659 ] = 8'h96;
  picture_data[ 1660 ] = 8'hE6;
  picture_data[ 1661 ] = 8'hB6;
  picture_data[ 1662 ] = 8'hDE;
  picture_data[ 1663 ] = 8'h55;
  picture_data[ 1664 ] = 8'hD6;
  picture_data[ 1665 ] = 8'h34;
  picture_data[ 1666 ] = 8'hDE;
  picture_data[ 1667 ] = 8'h74;
  picture_data[ 1668 ] = 8'hDE;
  picture_data[ 1669 ] = 8'h74;
  picture_data[ 1670 ] = 8'hD6;
  picture_data[ 1671 ] = 8'h33;
  picture_data[ 1672 ] = 8'h18;
  picture_data[ 1673 ] = 8'hA0;
  picture_data[ 1674 ] = 8'h18;
  picture_data[ 1675 ] = 8'hC0;
  picture_data[ 1676 ] = 8'h52;
  picture_data[ 1677 ] = 8'h87;
  picture_data[ 1678 ] = 8'h31;
  picture_data[ 1679 ] = 8'h83;
  picture_data[ 1680 ] = 8'h29;
  picture_data[ 1681 ] = 8'h42;
  picture_data[ 1682 ] = 8'h19;
  picture_data[ 1683 ] = 8'h01;
  picture_data[ 1684 ] = 8'h18;
  picture_data[ 1685 ] = 8'hE1;
  picture_data[ 1686 ] = 8'h19;
  picture_data[ 1687 ] = 8'h01;
  picture_data[ 1688 ] = 8'h10;
  picture_data[ 1689 ] = 8'hC1;
  picture_data[ 1690 ] = 8'h10;
  picture_data[ 1691 ] = 8'hE1;
  picture_data[ 1692 ] = 8'h18;
  picture_data[ 1693 ] = 8'hE2;
  picture_data[ 1694 ] = 8'h10;
  picture_data[ 1695 ] = 8'hE2;
  picture_data[ 1696 ] = 8'h21;
  picture_data[ 1697 ] = 8'h23;
  picture_data[ 1698 ] = 8'h19;
  picture_data[ 1699 ] = 8'h22;
  picture_data[ 1700 ] = 8'h29;
  picture_data[ 1701 ] = 8'h64;
  picture_data[ 1702 ] = 8'h21;
  picture_data[ 1703 ] = 8'h63;
  picture_data[ 1704 ] = 8'h29;
  picture_data[ 1705 ] = 8'hA5;
  picture_data[ 1706 ] = 8'h29;
  picture_data[ 1707 ] = 8'hC5;
  picture_data[ 1708 ] = 8'h19;
  picture_data[ 1709 ] = 8'h85;
  picture_data[ 1710 ] = 8'h19;
  picture_data[ 1711 ] = 8'h85;
  picture_data[ 1712 ] = 8'h21;
  picture_data[ 1713 ] = 8'hE7;
  picture_data[ 1714 ] = 8'h21;
  picture_data[ 1715 ] = 8'hA6;
  picture_data[ 1716 ] = 8'h19;
  picture_data[ 1717 ] = 8'h44;
  picture_data[ 1718 ] = 8'h19;
  picture_data[ 1719 ] = 8'h44;
  picture_data[ 1720 ] = 8'h09;
  picture_data[ 1721 ] = 8'h03;
  picture_data[ 1722 ] = 8'h11;
  picture_data[ 1723 ] = 8'h65;
  picture_data[ 1724 ] = 8'h11;
  picture_data[ 1725 ] = 8'h65;
  picture_data[ 1726 ] = 8'h11;
  picture_data[ 1727 ] = 8'h65;
  picture_data[ 1728 ] = 8'h11;
  picture_data[ 1729 ] = 8'h04;
  picture_data[ 1730 ] = 8'h11;
  picture_data[ 1731 ] = 8'h03;
  picture_data[ 1732 ] = 8'h08;
  picture_data[ 1733 ] = 8'hC2;
  picture_data[ 1734 ] = 8'h10;
  picture_data[ 1735 ] = 8'hE2;
  picture_data[ 1736 ] = 8'h21;
  picture_data[ 1737 ] = 8'h65;
  picture_data[ 1738 ] = 8'h21;
  picture_data[ 1739 ] = 8'h04;
  picture_data[ 1740 ] = 8'h18;
  picture_data[ 1741 ] = 8'h82;
  picture_data[ 1742 ] = 8'h31;
  picture_data[ 1743 ] = 8'h23;
  picture_data[ 1744 ] = 8'h39;
  picture_data[ 1745 ] = 8'h44;
  picture_data[ 1746 ] = 8'h49;
  picture_data[ 1747 ] = 8'h65;
  picture_data[ 1748 ] = 8'h59;
  picture_data[ 1749 ] = 8'h26;
  picture_data[ 1750 ] = 8'h60;
  picture_data[ 1751 ] = 8'hE5;
  picture_data[ 1752 ] = 8'h70;
  picture_data[ 1753 ] = 8'hE5;
  picture_data[ 1754 ] = 8'h68;
  picture_data[ 1755 ] = 8'hE5;
  picture_data[ 1756 ] = 8'h40;
  picture_data[ 1757 ] = 8'hC5;
  picture_data[ 1758 ] = 8'h20;
  picture_data[ 1759 ] = 8'hC8;
  picture_data[ 1760 ] = 8'h11;
  picture_data[ 1761 ] = 8'hB3;
  picture_data[ 1762 ] = 8'h2B;
  picture_data[ 1763 ] = 8'h5C;
  picture_data[ 1764 ] = 8'h2C;
  picture_data[ 1765 ] = 8'h5F;
  picture_data[ 1766 ] = 8'h23;
  picture_data[ 1767 ] = 8'hDA;
  picture_data[ 1768 ] = 8'h09;
  picture_data[ 1769 ] = 8'h8F;
  picture_data[ 1770 ] = 8'h19;
  picture_data[ 1771 ] = 8'h2B;
  picture_data[ 1772 ] = 8'h29;
  picture_data[ 1773 ] = 8'h69;
  picture_data[ 1774 ] = 8'h9C;
  picture_data[ 1775 ] = 8'hB3;
  picture_data[ 1776 ] = 8'hE6;
  picture_data[ 1777 ] = 8'hD9;
  picture_data[ 1778 ] = 8'hF7;
  picture_data[ 1779 ] = 8'h5A;
  picture_data[ 1780 ] = 8'hE6;
  picture_data[ 1781 ] = 8'hB8;
  picture_data[ 1782 ] = 8'hE6;
  picture_data[ 1783 ] = 8'h95;
  picture_data[ 1784 ] = 8'hCD;
  picture_data[ 1785 ] = 8'h6B;
  picture_data[ 1786 ] = 8'hB4;
  picture_data[ 1787 ] = 8'hA8;
  picture_data[ 1788 ] = 8'hBD;
  picture_data[ 1789 ] = 8'h2E;
  picture_data[ 1790 ] = 8'hEE;
  picture_data[ 1791 ] = 8'hF8;
  picture_data[ 1792 ] = 8'hFF;
  picture_data[ 1793 ] = 8'hFE;
  picture_data[ 1794 ] = 8'hC6;
  picture_data[ 1795 ] = 8'h17;
  picture_data[ 1796 ] = 8'hEE;
  picture_data[ 1797 ] = 8'hFB;
  picture_data[ 1798 ] = 8'hFF;
  picture_data[ 1799 ] = 8'hDE;
  picture_data[ 1800 ] = 8'hFF;
  picture_data[ 1801 ] = 8'hBC;
  picture_data[ 1802 ] = 8'hFF;
  picture_data[ 1803 ] = 8'hBB;
  picture_data[ 1804 ] = 8'hEF;
  picture_data[ 1805 ] = 8'h39;
  picture_data[ 1806 ] = 8'hE6;
  picture_data[ 1807 ] = 8'hF8;
  picture_data[ 1808 ] = 8'hE6;
  picture_data[ 1809 ] = 8'hD8;
  picture_data[ 1810 ] = 8'hE6;
  picture_data[ 1811 ] = 8'h96;
  picture_data[ 1812 ] = 8'hE6;
  picture_data[ 1813 ] = 8'h96;
  picture_data[ 1814 ] = 8'hDE;
  picture_data[ 1815 ] = 8'h95;
  picture_data[ 1816 ] = 8'hE6;
  picture_data[ 1817 ] = 8'h95;
  picture_data[ 1818 ] = 8'hDE;
  picture_data[ 1819 ] = 8'h74;
  picture_data[ 1820 ] = 8'hDE;
  picture_data[ 1821 ] = 8'h74;
  picture_data[ 1822 ] = 8'hD6;
  picture_data[ 1823 ] = 8'h53;
  picture_data[ 1824 ] = 8'h18;
  picture_data[ 1825 ] = 8'hC1;
  picture_data[ 1826 ] = 8'h18;
  picture_data[ 1827 ] = 8'hC0;
  picture_data[ 1828 ] = 8'h10;
  picture_data[ 1829 ] = 8'h80;
  picture_data[ 1830 ] = 8'h10;
  picture_data[ 1831 ] = 8'hA0;
  picture_data[ 1832 ] = 8'h10;
  picture_data[ 1833 ] = 8'hA0;
  picture_data[ 1834 ] = 8'h19;
  picture_data[ 1835 ] = 8'h02;
  picture_data[ 1836 ] = 8'h10;
  picture_data[ 1837 ] = 8'hA0;
  picture_data[ 1838 ] = 8'h18;
  picture_data[ 1839 ] = 8'hE2;
  picture_data[ 1840 ] = 8'h10;
  picture_data[ 1841 ] = 8'hC1;
  picture_data[ 1842 ] = 8'h19;
  picture_data[ 1843 ] = 8'h02;
  picture_data[ 1844 ] = 8'h10;
  picture_data[ 1845 ] = 8'hE2;
  picture_data[ 1846 ] = 8'h08;
  picture_data[ 1847 ] = 8'hA1;
  picture_data[ 1848 ] = 8'h18;
  picture_data[ 1849 ] = 8'hE2;
  picture_data[ 1850 ] = 8'h21;
  picture_data[ 1851 ] = 8'h22;
  picture_data[ 1852 ] = 8'h21;
  picture_data[ 1853 ] = 8'h23;
  picture_data[ 1854 ] = 8'h19;
  picture_data[ 1855 ] = 8'h02;
  picture_data[ 1856 ] = 8'h19;
  picture_data[ 1857 ] = 8'h43;
  picture_data[ 1858 ] = 8'h11;
  picture_data[ 1859 ] = 8'h43;
  picture_data[ 1860 ] = 8'h21;
  picture_data[ 1861 ] = 8'hE6;
  picture_data[ 1862 ] = 8'h22;
  picture_data[ 1863 ] = 8'h07;
  picture_data[ 1864 ] = 8'h11;
  picture_data[ 1865 ] = 8'h44;
  picture_data[ 1866 ] = 8'h11;
  picture_data[ 1867 ] = 8'h24;
  picture_data[ 1868 ] = 8'h11;
  picture_data[ 1869 ] = 8'h04;
  picture_data[ 1870 ] = 8'h08;
  picture_data[ 1871 ] = 8'hC2;
  picture_data[ 1872 ] = 8'h09;
  picture_data[ 1873 ] = 8'h24;
  picture_data[ 1874 ] = 8'h09;
  picture_data[ 1875 ] = 8'h44;
  picture_data[ 1876 ] = 8'h11;
  picture_data[ 1877 ] = 8'h65;
  picture_data[ 1878 ] = 8'h19;
  picture_data[ 1879 ] = 8'hA6;
  picture_data[ 1880 ] = 8'h19;
  picture_data[ 1881 ] = 8'h65;
  picture_data[ 1882 ] = 8'h11;
  picture_data[ 1883 ] = 8'h24;
  picture_data[ 1884 ] = 8'h11;
  picture_data[ 1885 ] = 8'h23;
  picture_data[ 1886 ] = 8'h19;
  picture_data[ 1887 ] = 8'h44;
  picture_data[ 1888 ] = 8'h11;
  picture_data[ 1889 ] = 8'h24;
  picture_data[ 1890 ] = 8'h10;
  picture_data[ 1891 ] = 8'hC3;
  picture_data[ 1892 ] = 8'h18;
  picture_data[ 1893 ] = 8'h82;
  picture_data[ 1894 ] = 8'h28;
  picture_data[ 1895 ] = 8'hE4;
  picture_data[ 1896 ] = 8'h31;
  picture_data[ 1897 ] = 8'h24;
  picture_data[ 1898 ] = 8'h31;
  picture_data[ 1899 ] = 8'h44;
  picture_data[ 1900 ] = 8'h39;
  picture_data[ 1901 ] = 8'h04;
  picture_data[ 1902 ] = 8'h41;
  picture_data[ 1903 ] = 8'h05;
  picture_data[ 1904 ] = 8'h49;
  picture_data[ 1905 ] = 8'h05;
  picture_data[ 1906 ] = 8'h49;
  picture_data[ 1907 ] = 8'h46;
  picture_data[ 1908 ] = 8'h29;
  picture_data[ 1909 ] = 8'h26;
  picture_data[ 1910 ] = 8'h19;
  picture_data[ 1911 ] = 8'h49;
  picture_data[ 1912 ] = 8'h11;
  picture_data[ 1913 ] = 8'h70;
  picture_data[ 1914 ] = 8'h2A;
  picture_data[ 1915 ] = 8'hB8;
  picture_data[ 1916 ] = 8'h44;
  picture_data[ 1917 ] = 8'h3C;
  picture_data[ 1918 ] = 8'h3B;
  picture_data[ 1919 ] = 8'hD8;
  picture_data[ 1920 ] = 8'h7C;
  picture_data[ 1921 ] = 8'h97;
  picture_data[ 1922 ] = 8'h6B;
  picture_data[ 1923 ] = 8'h70;
  picture_data[ 1924 ] = 8'h5B;
  picture_data[ 1925 ] = 8'h0D;
  picture_data[ 1926 ] = 8'h9C;
  picture_data[ 1927 ] = 8'hF3;
  picture_data[ 1928 ] = 8'hC6;
  picture_data[ 1929 ] = 8'h37;
  picture_data[ 1930 ] = 8'hFF;
  picture_data[ 1931 ] = 8'hFE;
  picture_data[ 1932 ] = 8'hFF;
  picture_data[ 1933 ] = 8'hFE;
  picture_data[ 1934 ] = 8'hFF;
  picture_data[ 1935 ] = 8'hFC;
  picture_data[ 1936 ] = 8'hDE;
  picture_data[ 1937 ] = 8'h31;
  picture_data[ 1938 ] = 8'hBD;
  picture_data[ 1939 ] = 8'h2C;
  picture_data[ 1940 ] = 8'hE6;
  picture_data[ 1941 ] = 8'h95;
  picture_data[ 1942 ] = 8'hD6;
  picture_data[ 1943 ] = 8'h96;
  picture_data[ 1944 ] = 8'hFF;
  picture_data[ 1945 ] = 8'hFD;
  picture_data[ 1946 ] = 8'hBD;
  picture_data[ 1947 ] = 8'hD5;
  picture_data[ 1948 ] = 8'hEF;
  picture_data[ 1949 ] = 8'h1A;
  picture_data[ 1950 ] = 8'hFF;
  picture_data[ 1951 ] = 8'hFD;
  picture_data[ 1952 ] = 8'hFF;
  picture_data[ 1953 ] = 8'hDC;
  picture_data[ 1954 ] = 8'hF7;
  picture_data[ 1955 ] = 8'h9B;
  picture_data[ 1956 ] = 8'hEF;
  picture_data[ 1957 ] = 8'h39;
  picture_data[ 1958 ] = 8'hF7;
  picture_data[ 1959 ] = 8'h9A;
  picture_data[ 1960 ] = 8'hF7;
  picture_data[ 1961 ] = 8'h59;
  picture_data[ 1962 ] = 8'hF7;
  picture_data[ 1963 ] = 8'h39;
  picture_data[ 1964 ] = 8'hF7;
  picture_data[ 1965 ] = 8'h18;
  picture_data[ 1966 ] = 8'hEE;
  picture_data[ 1967 ] = 8'hD7;
  picture_data[ 1968 ] = 8'hEE;
  picture_data[ 1969 ] = 8'hD6;
  picture_data[ 1970 ] = 8'hE6;
  picture_data[ 1971 ] = 8'h95;
  picture_data[ 1972 ] = 8'hE6;
  picture_data[ 1973 ] = 8'h95;
  picture_data[ 1974 ] = 8'hDE;
  picture_data[ 1975 ] = 8'h33;
  picture_data[ 1976 ] = 8'h10;
  picture_data[ 1977 ] = 8'hA1;
  picture_data[ 1978 ] = 8'h10;
  picture_data[ 1979 ] = 8'hC1;
  picture_data[ 1980 ] = 8'h10;
  picture_data[ 1981 ] = 8'hC1;
  picture_data[ 1982 ] = 8'h08;
  picture_data[ 1983 ] = 8'hA1;
  picture_data[ 1984 ] = 8'h10;
  picture_data[ 1985 ] = 8'hE2;
  picture_data[ 1986 ] = 8'h19;
  picture_data[ 1987 ] = 8'h02;
  picture_data[ 1988 ] = 8'h21;
  picture_data[ 1989 ] = 8'h43;
  picture_data[ 1990 ] = 8'h10;
  picture_data[ 1991 ] = 8'hA1;
  picture_data[ 1992 ] = 8'h10;
  picture_data[ 1993 ] = 8'hA1;
  picture_data[ 1994 ] = 8'h10;
  picture_data[ 1995 ] = 8'hA1;
  picture_data[ 1996 ] = 8'h10;
  picture_data[ 1997 ] = 8'hC2;
  picture_data[ 1998 ] = 8'h10;
  picture_data[ 1999 ] = 8'hE2;
  picture_data[ 2000 ] = 8'h21;
  picture_data[ 2001 ] = 8'h23;
  picture_data[ 2002 ] = 8'h29;
  picture_data[ 2003 ] = 8'h43;
  picture_data[ 2004 ] = 8'h21;
  picture_data[ 2005 ] = 8'h02;
  picture_data[ 2006 ] = 8'h29;
  picture_data[ 2007 ] = 8'h42;
  picture_data[ 2008 ] = 8'h21;
  picture_data[ 2009 ] = 8'h43;
  picture_data[ 2010 ] = 8'h21;
  picture_data[ 2011 ] = 8'hA4;
  picture_data[ 2012 ] = 8'h32;
  picture_data[ 2013 ] = 8'h68;
  picture_data[ 2014 ] = 8'h21;
  picture_data[ 2015 ] = 8'hE6;
  picture_data[ 2016 ] = 8'h08;
  picture_data[ 2017 ] = 8'hE3;
  picture_data[ 2018 ] = 8'h09;
  picture_data[ 2019 ] = 8'h04;
  picture_data[ 2020 ] = 8'h10;
  picture_data[ 2021 ] = 8'hE3;
  picture_data[ 2022 ] = 8'h08;
  picture_data[ 2023 ] = 8'hA2;
  picture_data[ 2024 ] = 8'h09;
  picture_data[ 2025 ] = 8'h23;
  picture_data[ 2026 ] = 8'h09;
  picture_data[ 2027 ] = 8'h23;
  picture_data[ 2028 ] = 8'h09;
  picture_data[ 2029 ] = 8'h44;
  picture_data[ 2030 ] = 8'h11;
  picture_data[ 2031 ] = 8'h65;
  picture_data[ 2032 ] = 8'h11;
  picture_data[ 2033 ] = 8'h24;
  picture_data[ 2034 ] = 8'h11;
  picture_data[ 2035 ] = 8'h24;
  picture_data[ 2036 ] = 8'h11;
  picture_data[ 2037 ] = 8'h44;
  picture_data[ 2038 ] = 8'h19;
  picture_data[ 2039 ] = 8'h44;
  picture_data[ 2040 ] = 8'h32;
  picture_data[ 2041 ] = 8'h08;
  picture_data[ 2042 ] = 8'h21;
  picture_data[ 2043 ] = 8'h45;
  picture_data[ 2044 ] = 8'h21;
  picture_data[ 2045 ] = 8'h04;
  picture_data[ 2046 ] = 8'h20;
  picture_data[ 2047 ] = 8'hE3;
  picture_data[ 2048 ] = 8'h18;
  picture_data[ 2049 ] = 8'hE2;
  picture_data[ 2050 ] = 8'h18;
  picture_data[ 2051 ] = 8'hC1;
  picture_data[ 2052 ] = 8'h29;
  picture_data[ 2053 ] = 8'h03;
  picture_data[ 2054 ] = 8'h31;
  picture_data[ 2055 ] = 8'h45;
  picture_data[ 2056 ] = 8'h39;
  picture_data[ 2057 ] = 8'h46;
  picture_data[ 2058 ] = 8'h20;
  picture_data[ 2059 ] = 8'hE4;
  picture_data[ 2060 ] = 8'h29;
  picture_data[ 2061 ] = 8'h66;
  picture_data[ 2062 ] = 8'h21;
  picture_data[ 2063 ] = 8'h68;
  picture_data[ 2064 ] = 8'h08;
  picture_data[ 2065 ] = 8'hCA;
  picture_data[ 2066 ] = 8'h4B;
  picture_data[ 2067 ] = 8'h14;
  picture_data[ 2068 ] = 8'h64;
  picture_data[ 2069 ] = 8'h37;
  picture_data[ 2070 ] = 8'h9D;
  picture_data[ 2071 ] = 8'hBC;
  picture_data[ 2072 ] = 8'hFF;
  picture_data[ 2073 ] = 8'hFF;
  picture_data[ 2074 ] = 8'hFF;
  picture_data[ 2075 ] = 8'hDF;
  picture_data[ 2076 ] = 8'hF7;
  picture_data[ 2077 ] = 8'h9E;
  picture_data[ 2078 ] = 8'hD6;
  picture_data[ 2079 ] = 8'hBA;
  picture_data[ 2080 ] = 8'hB5;
  picture_data[ 2081 ] = 8'h95;
  picture_data[ 2082 ] = 8'h7B;
  picture_data[ 2083 ] = 8'hEE;
  picture_data[ 2084 ] = 8'hA5;
  picture_data[ 2085 ] = 8'h13;
  picture_data[ 2086 ] = 8'hFF;
  picture_data[ 2087 ] = 8'hFD;
  picture_data[ 2088 ] = 8'hBD;
  picture_data[ 2089 ] = 8'h50;
  picture_data[ 2090 ] = 8'hFF;
  picture_data[ 2091 ] = 8'h57;
  picture_data[ 2092 ] = 8'hEE;
  picture_data[ 2093 ] = 8'hF8;
  picture_data[ 2094 ] = 8'hCE;
  picture_data[ 2095 ] = 8'h76;
  picture_data[ 2096 ] = 8'hEF;
  picture_data[ 2097 ] = 8'h5B;
  picture_data[ 2098 ] = 8'hBD;
  picture_data[ 2099 ] = 8'hB4;
  picture_data[ 2100 ] = 8'hD6;
  picture_data[ 2101 ] = 8'h56;
  picture_data[ 2102 ] = 8'hEF;
  picture_data[ 2103 ] = 8'h19;
  picture_data[ 2104 ] = 8'hD6;
  picture_data[ 2105 ] = 8'h77;
  picture_data[ 2106 ] = 8'hF7;
  picture_data[ 2107 ] = 8'h5A;
  picture_data[ 2108 ] = 8'hF7;
  picture_data[ 2109 ] = 8'h7A;
  picture_data[ 2110 ] = 8'hEF;
  picture_data[ 2111 ] = 8'h19;
  picture_data[ 2112 ] = 8'hE6;
  picture_data[ 2113 ] = 8'hB7;
  picture_data[ 2114 ] = 8'hE6;
  picture_data[ 2115 ] = 8'h96;
  picture_data[ 2116 ] = 8'hDE;
  picture_data[ 2117 ] = 8'h55;
  picture_data[ 2118 ] = 8'hD6;
  picture_data[ 2119 ] = 8'h34;
  picture_data[ 2120 ] = 8'hCD;
  picture_data[ 2121 ] = 8'hB2;
  picture_data[ 2122 ] = 8'hDE;
  picture_data[ 2123 ] = 8'h34;
  picture_data[ 2124 ] = 8'hEE;
  picture_data[ 2125 ] = 8'hD6;
  picture_data[ 2126 ] = 8'hDE;
  picture_data[ 2127 ] = 8'h34;
  picture_data[ 2128 ] = 8'h08;
  picture_data[ 2129 ] = 8'h61;
  picture_data[ 2130 ] = 8'h10;
  picture_data[ 2131 ] = 8'hC2;
  picture_data[ 2132 ] = 8'h08;
  picture_data[ 2133 ] = 8'hA2;
  picture_data[ 2134 ] = 8'h08;
  picture_data[ 2135 ] = 8'hC2;
  picture_data[ 2136 ] = 8'h08;
  picture_data[ 2137 ] = 8'hA1;
  picture_data[ 2138 ] = 8'h10;
  picture_data[ 2139 ] = 8'hE2;
  picture_data[ 2140 ] = 8'h18;
  picture_data[ 2141 ] = 8'hE3;
  picture_data[ 2142 ] = 8'h10;
  picture_data[ 2143 ] = 8'hC2;
  picture_data[ 2144 ] = 8'h21;
  picture_data[ 2145 ] = 8'h03;
  picture_data[ 2146 ] = 8'h10;
  picture_data[ 2147 ] = 8'hA1;
  picture_data[ 2148 ] = 8'h19;
  picture_data[ 2149 ] = 8'h02;
  picture_data[ 2150 ] = 8'h19;
  picture_data[ 2151 ] = 8'h22;
  picture_data[ 2152 ] = 8'h10;
  picture_data[ 2153 ] = 8'hC1;
  picture_data[ 2154 ] = 8'h29;
  picture_data[ 2155 ] = 8'h63;
  picture_data[ 2156 ] = 8'h29;
  picture_data[ 2157 ] = 8'h22;
  picture_data[ 2158 ] = 8'h20;
  picture_data[ 2159 ] = 8'hE1;
  picture_data[ 2160 ] = 8'h21;
  picture_data[ 2161 ] = 8'h42;
  picture_data[ 2162 ] = 8'h29;
  picture_data[ 2163 ] = 8'hE5;
  picture_data[ 2164 ] = 8'h42;
  picture_data[ 2165 ] = 8'hA8;
  picture_data[ 2166 ] = 8'h09;
  picture_data[ 2167 ] = 8'h43;
  picture_data[ 2168 ] = 8'h00;
  picture_data[ 2169 ] = 8'hC2;
  picture_data[ 2170 ] = 8'h08;
  picture_data[ 2171 ] = 8'hC2;
  picture_data[ 2172 ] = 8'h08;
  picture_data[ 2173 ] = 8'hA1;
  picture_data[ 2174 ] = 8'h11;
  picture_data[ 2175 ] = 8'h03;
  picture_data[ 2176 ] = 8'h11;
  picture_data[ 2177 ] = 8'h23;
  picture_data[ 2178 ] = 8'h09;
  picture_data[ 2179 ] = 8'h23;
  picture_data[ 2180 ] = 8'h09;
  picture_data[ 2181 ] = 8'h24;
  picture_data[ 2182 ] = 8'h11;
  picture_data[ 2183 ] = 8'h65;
  picture_data[ 2184 ] = 8'h11;
  picture_data[ 2185 ] = 8'h24;
  picture_data[ 2186 ] = 8'h08;
  picture_data[ 2187 ] = 8'hE3;
  picture_data[ 2188 ] = 8'h11;
  picture_data[ 2189 ] = 8'h02;
  picture_data[ 2190 ] = 8'h21;
  picture_data[ 2191 ] = 8'h64;
  picture_data[ 2192 ] = 8'h19;
  picture_data[ 2193 ] = 8'h24;
  picture_data[ 2194 ] = 8'h29;
  picture_data[ 2195 ] = 8'hA6;
  picture_data[ 2196 ] = 8'h29;
  picture_data[ 2197 ] = 8'h85;
  picture_data[ 2198 ] = 8'h19;
  picture_data[ 2199 ] = 8'h43;
  picture_data[ 2200 ] = 8'h29;
  picture_data[ 2201 ] = 8'hC3;
  picture_data[ 2202 ] = 8'h29;
  picture_data[ 2203 ] = 8'h83;
  picture_data[ 2204 ] = 8'h29;
  picture_data[ 2205 ] = 8'h23;
  picture_data[ 2206 ] = 8'h28;
  picture_data[ 2207 ] = 8'hE3;
  picture_data[ 2208 ] = 8'h20;
  picture_data[ 2209 ] = 8'hA4;
  picture_data[ 2210 ] = 8'h20;
  picture_data[ 2211 ] = 8'hC4;
  picture_data[ 2212 ] = 8'h20;
  picture_data[ 2213 ] = 8'hA2;
  picture_data[ 2214 ] = 8'h39;
  picture_data[ 2215 ] = 8'hC6;
  picture_data[ 2216 ] = 8'h7B;
  picture_data[ 2217 ] = 8'h8E;
  picture_data[ 2218 ] = 8'h6B;
  picture_data[ 2219 ] = 8'h6E;
  picture_data[ 2220 ] = 8'h9C;
  picture_data[ 2221 ] = 8'hF3;
  picture_data[ 2222 ] = 8'hF7;
  picture_data[ 2223 ] = 8'h9D;
  picture_data[ 2224 ] = 8'hFF;
  picture_data[ 2225 ] = 8'hBF;
  picture_data[ 2226 ] = 8'hFF;
  picture_data[ 2227 ] = 8'hBF;
  picture_data[ 2228 ] = 8'hFF;
  picture_data[ 2229 ] = 8'hFF;
  picture_data[ 2230 ] = 8'hB5;
  picture_data[ 2231 ] = 8'h97;
  picture_data[ 2232 ] = 8'h5A;
  picture_data[ 2233 ] = 8'hAC;
  picture_data[ 2234 ] = 8'h4A;
  picture_data[ 2235 ] = 8'h29;
  picture_data[ 2236 ] = 8'h8C;
  picture_data[ 2237 ] = 8'h50;
  picture_data[ 2238 ] = 8'hEE;
  picture_data[ 2239 ] = 8'hFA;
  picture_data[ 2240 ] = 8'h9C;
  picture_data[ 2241 ] = 8'h2E;
  picture_data[ 2242 ] = 8'hB5;
  picture_data[ 2243 ] = 8'h11;
  picture_data[ 2244 ] = 8'h94;
  picture_data[ 2245 ] = 8'h4E;
  picture_data[ 2246 ] = 8'h6B;
  picture_data[ 2247 ] = 8'h2A;
  picture_data[ 2248 ] = 8'h52;
  picture_data[ 2249 ] = 8'h67;
  picture_data[ 2250 ] = 8'h5A;
  picture_data[ 2251 ] = 8'h88;
  picture_data[ 2252 ] = 8'h4A;
  picture_data[ 2253 ] = 8'h25;
  picture_data[ 2254 ] = 8'h49;
  picture_data[ 2255 ] = 8'hE4;
  picture_data[ 2256 ] = 8'h6A;
  picture_data[ 2257 ] = 8'hA7;
  picture_data[ 2258 ] = 8'hA4;
  picture_data[ 2259 ] = 8'h6E;
  picture_data[ 2260 ] = 8'hE6;
  picture_data[ 2261 ] = 8'h76;
  picture_data[ 2262 ] = 8'hE6;
  picture_data[ 2263 ] = 8'h96;
  picture_data[ 2264 ] = 8'h9C;
  picture_data[ 2265 ] = 8'h2D;
  picture_data[ 2266 ] = 8'hA4;
  picture_data[ 2267 ] = 8'h4D;
  picture_data[ 2268 ] = 8'hAC;
  picture_data[ 2269 ] = 8'hCF;
  picture_data[ 2270 ] = 8'hA4;
  picture_data[ 2271 ] = 8'hAE;
  picture_data[ 2272 ] = 8'hAC;
  picture_data[ 2273 ] = 8'hAE;
  picture_data[ 2274 ] = 8'hCD;
  picture_data[ 2275 ] = 8'hD2;
  picture_data[ 2276 ] = 8'hF6;
  picture_data[ 2277 ] = 8'hF7;
  picture_data[ 2278 ] = 8'hDE;
  picture_data[ 2279 ] = 8'h75;
  picture_data[ 2280 ] = 8'h10;
  picture_data[ 2281 ] = 8'hE3;
  picture_data[ 2282 ] = 8'h08;
  picture_data[ 2283 ] = 8'h82;
  picture_data[ 2284 ] = 8'h10;
  picture_data[ 2285 ] = 8'hE3;
  picture_data[ 2286 ] = 8'h11;
  picture_data[ 2287 ] = 8'h04;
  picture_data[ 2288 ] = 8'h10;
  picture_data[ 2289 ] = 8'hE3;
  picture_data[ 2290 ] = 8'h08;
  picture_data[ 2291 ] = 8'hC2;
  picture_data[ 2292 ] = 8'h10;
  picture_data[ 2293 ] = 8'hC2;
  picture_data[ 2294 ] = 8'h18;
  picture_data[ 2295 ] = 8'hE2;
  picture_data[ 2296 ] = 8'h18;
  picture_data[ 2297 ] = 8'hC2;
  picture_data[ 2298 ] = 8'h18;
  picture_data[ 2299 ] = 8'hE2;
  picture_data[ 2300 ] = 8'h19;
  picture_data[ 2301 ] = 8'h03;
  picture_data[ 2302 ] = 8'h21;
  picture_data[ 2303 ] = 8'h23;
  picture_data[ 2304 ] = 8'h29;
  picture_data[ 2305 ] = 8'h22;
  picture_data[ 2306 ] = 8'h39;
  picture_data[ 2307 ] = 8'h82;
  picture_data[ 2308 ] = 8'h41;
  picture_data[ 2309 ] = 8'h81;
  picture_data[ 2310 ] = 8'h7B;
  picture_data[ 2311 ] = 8'h68;
  picture_data[ 2312 ] = 8'h83;
  picture_data[ 2313 ] = 8'hC9;
  picture_data[ 2314 ] = 8'h62;
  picture_data[ 2315 ] = 8'hE6;
  picture_data[ 2316 ] = 8'h52;
  picture_data[ 2317 ] = 8'hE8;
  picture_data[ 2318 ] = 8'h08;
  picture_data[ 2319 ] = 8'hE2;
  picture_data[ 2320 ] = 8'h08;
  picture_data[ 2321 ] = 8'hC2;
  picture_data[ 2322 ] = 8'h10;
  picture_data[ 2323 ] = 8'hE3;
  picture_data[ 2324 ] = 8'h10;
  picture_data[ 2325 ] = 8'hE2;
  picture_data[ 2326 ] = 8'h11;
  picture_data[ 2327 ] = 8'h02;
  picture_data[ 2328 ] = 8'h11;
  picture_data[ 2329 ] = 8'h03;
  picture_data[ 2330 ] = 8'h11;
  picture_data[ 2331 ] = 8'h64;
  picture_data[ 2332 ] = 8'h11;
  picture_data[ 2333 ] = 8'h64;
  picture_data[ 2334 ] = 8'h11;
  picture_data[ 2335 ] = 8'h65;
  picture_data[ 2336 ] = 8'h19;
  picture_data[ 2337 ] = 8'h65;
  picture_data[ 2338 ] = 8'h08;
  picture_data[ 2339 ] = 8'hE3;
  picture_data[ 2340 ] = 8'h08;
  picture_data[ 2341 ] = 8'hC2;
  picture_data[ 2342 ] = 8'h19;
  picture_data[ 2343 ] = 8'h44;
  picture_data[ 2344 ] = 8'h19;
  picture_data[ 2345 ] = 8'h45;
  picture_data[ 2346 ] = 8'h19;
  picture_data[ 2347 ] = 8'h44;
  picture_data[ 2348 ] = 8'h11;
  picture_data[ 2349 ] = 8'h22;
  picture_data[ 2350 ] = 8'h29;
  picture_data[ 2351 ] = 8'hE5;
  picture_data[ 2352 ] = 8'h21;
  picture_data[ 2353 ] = 8'hA3;
  picture_data[ 2354 ] = 8'h21;
  picture_data[ 2355 ] = 8'h42;
  picture_data[ 2356 ] = 8'h29;
  picture_data[ 2357 ] = 8'h43;
  picture_data[ 2358 ] = 8'h39;
  picture_data[ 2359 ] = 8'h65;
  picture_data[ 2360 ] = 8'h41;
  picture_data[ 2361 ] = 8'hC7;
  picture_data[ 2362 ] = 8'h41;
  picture_data[ 2363 ] = 8'hA6;
  picture_data[ 2364 ] = 8'h6A;
  picture_data[ 2365 ] = 8'hEA;
  picture_data[ 2366 ] = 8'hA4;
  picture_data[ 2367 ] = 8'h8F;
  picture_data[ 2368 ] = 8'hDE;
  picture_data[ 2369 ] = 8'h77;
  picture_data[ 2370 ] = 8'hC5;
  picture_data[ 2371 ] = 8'h93;
  picture_data[ 2372 ] = 8'hC5;
  picture_data[ 2373 ] = 8'h72;
  picture_data[ 2374 ] = 8'hF7;
  picture_data[ 2375 ] = 8'h3A;
  picture_data[ 2376 ] = 8'hFF;
  picture_data[ 2377 ] = 8'h7D;
  picture_data[ 2378 ] = 8'hD5;
  picture_data[ 2379 ] = 8'hF9;
  picture_data[ 2380 ] = 8'h83;
  picture_data[ 2381 ] = 8'hB0;
  picture_data[ 2382 ] = 8'h4A;
  picture_data[ 2383 ] = 8'h2A;
  picture_data[ 2384 ] = 8'h6A;
  picture_data[ 2385 ] = 8'hEE;
  picture_data[ 2386 ] = 8'h52;
  picture_data[ 2387 ] = 8'h4B;
  picture_data[ 2388 ] = 8'h73;
  picture_data[ 2389 ] = 8'h8D;
  picture_data[ 2390 ] = 8'hB5;
  picture_data[ 2391 ] = 8'h54;
  picture_data[ 2392 ] = 8'h8B;
  picture_data[ 2393 ] = 8'hAE;
  picture_data[ 2394 ] = 8'h39;
  picture_data[ 2395 ] = 8'h24;
  picture_data[ 2396 ] = 8'h29;
  picture_data[ 2397 ] = 8'h02;
  picture_data[ 2398 ] = 8'h41;
  picture_data[ 2399 ] = 8'hC4;
  picture_data[ 2400 ] = 8'h49;
  picture_data[ 2401 ] = 8'hE5;
  picture_data[ 2402 ] = 8'h52;
  picture_data[ 2403 ] = 8'h05;
  picture_data[ 2404 ] = 8'h49;
  picture_data[ 2405 ] = 8'hE4;
  picture_data[ 2406 ] = 8'h41;
  picture_data[ 2407 ] = 8'h62;
  picture_data[ 2408 ] = 8'h51;
  picture_data[ 2409 ] = 8'h82;
  picture_data[ 2410 ] = 8'h61;
  picture_data[ 2411 ] = 8'hC4;
  picture_data[ 2412 ] = 8'h72;
  picture_data[ 2413 ] = 8'h25;
  picture_data[ 2414 ] = 8'h6A;
  picture_data[ 2415 ] = 8'h25;
  picture_data[ 2416 ] = 8'hAC;
  picture_data[ 2417 ] = 8'h8E;
  picture_data[ 2418 ] = 8'hBC;
  picture_data[ 2419 ] = 8'hF0;
  picture_data[ 2420 ] = 8'hB4;
  picture_data[ 2421 ] = 8'hEF;
  picture_data[ 2422 ] = 8'hB5;
  picture_data[ 2423 ] = 8'h10;
  picture_data[ 2424 ] = 8'hB4;
  picture_data[ 2425 ] = 8'hEF;
  picture_data[ 2426 ] = 8'hCD;
  picture_data[ 2427 ] = 8'hB2;
  picture_data[ 2428 ] = 8'hEE;
  picture_data[ 2429 ] = 8'hF7;
  picture_data[ 2430 ] = 8'hE6;
  picture_data[ 2431 ] = 8'h96;
  picture_data[ 2432 ] = 8'h08;
  picture_data[ 2433 ] = 8'hC2;
  picture_data[ 2434 ] = 8'h08;
  picture_data[ 2435 ] = 8'hC2;
  picture_data[ 2436 ] = 8'h00;
  picture_data[ 2437 ] = 8'hA2;
  picture_data[ 2438 ] = 8'h00;
  picture_data[ 2439 ] = 8'h61;
  picture_data[ 2440 ] = 8'h08;
  picture_data[ 2441 ] = 8'hA2;
  picture_data[ 2442 ] = 8'h10;
  picture_data[ 2443 ] = 8'hC3;
  picture_data[ 2444 ] = 8'h10;
  picture_data[ 2445 ] = 8'hE2;
  picture_data[ 2446 ] = 8'h10;
  picture_data[ 2447 ] = 8'hC2;
  picture_data[ 2448 ] = 8'h19;
  picture_data[ 2449 ] = 8'h02;
  picture_data[ 2450 ] = 8'h21;
  picture_data[ 2451 ] = 8'h44;
  picture_data[ 2452 ] = 8'h31;
  picture_data[ 2453 ] = 8'h86;
  picture_data[ 2454 ] = 8'h20;
  picture_data[ 2455 ] = 8'hC2;
  picture_data[ 2456 ] = 8'h31;
  picture_data[ 2457 ] = 8'h22;
  picture_data[ 2458 ] = 8'h31;
  picture_data[ 2459 ] = 8'h00;
  picture_data[ 2460 ] = 8'h6A;
  picture_data[ 2461 ] = 8'h81;
  picture_data[ 2462 ] = 8'hE6;
  picture_data[ 2463 ] = 8'h0D;
  picture_data[ 2464 ] = 8'hEE;
  picture_data[ 2465 ] = 8'h4D;
  picture_data[ 2466 ] = 8'hDD;
  picture_data[ 2467 ] = 8'hCD;
  picture_data[ 2468 ] = 8'h5A;
  picture_data[ 2469 ] = 8'h45;
  picture_data[ 2470 ] = 8'h18;
  picture_data[ 2471 ] = 8'hA1;
  picture_data[ 2472 ] = 8'h10;
  picture_data[ 2473 ] = 8'hC2;
  picture_data[ 2474 ] = 8'h08;
  picture_data[ 2475 ] = 8'hA2;
  picture_data[ 2476 ] = 8'h10;
  picture_data[ 2477 ] = 8'hE3;
  picture_data[ 2478 ] = 8'h11;
  picture_data[ 2479 ] = 8'h02;
  picture_data[ 2480 ] = 8'h19;
  picture_data[ 2481 ] = 8'h43;
  picture_data[ 2482 ] = 8'h19;
  picture_data[ 2483 ] = 8'h43;
  picture_data[ 2484 ] = 8'h11;
  picture_data[ 2485 ] = 8'h03;
  picture_data[ 2486 ] = 8'h19;
  picture_data[ 2487 ] = 8'h45;
  picture_data[ 2488 ] = 8'h29;
  picture_data[ 2489 ] = 8'hC8;
  picture_data[ 2490 ] = 8'h19;
  picture_data[ 2491 ] = 8'h46;
  picture_data[ 2492 ] = 8'h11;
  picture_data[ 2493 ] = 8'h44;
  picture_data[ 2494 ] = 8'h21;
  picture_data[ 2495 ] = 8'h85;
  picture_data[ 2496 ] = 8'h19;
  picture_data[ 2497 ] = 8'h65;
  picture_data[ 2498 ] = 8'h21;
  picture_data[ 2499 ] = 8'h65;
  picture_data[ 2500 ] = 8'h21;
  picture_data[ 2501 ] = 8'h64;
  picture_data[ 2502 ] = 8'h29;
  picture_data[ 2503 ] = 8'h84;
  picture_data[ 2504 ] = 8'h29;
  picture_data[ 2505 ] = 8'h63;
  picture_data[ 2506 ] = 8'h29;
  picture_data[ 2507 ] = 8'h43;
  picture_data[ 2508 ] = 8'h20;
  picture_data[ 2509 ] = 8'hC2;
  picture_data[ 2510 ] = 8'h31;
  picture_data[ 2511 ] = 8'h24;
  picture_data[ 2512 ] = 8'h5A;
  picture_data[ 2513 ] = 8'h28;
  picture_data[ 2514 ] = 8'h83;
  picture_data[ 2515 ] = 8'h6C;
  picture_data[ 2516 ] = 8'hCD;
  picture_data[ 2517 ] = 8'hB4;
  picture_data[ 2518 ] = 8'hC5;
  picture_data[ 2519 ] = 8'h93;
  picture_data[ 2520 ] = 8'hCD;
  picture_data[ 2521 ] = 8'hD4;
  picture_data[ 2522 ] = 8'hD6;
  picture_data[ 2523 ] = 8'h36;
  picture_data[ 2524 ] = 8'hD6;
  picture_data[ 2525 ] = 8'h16;
  picture_data[ 2526 ] = 8'h83;
  picture_data[ 2527 ] = 8'h8D;
  picture_data[ 2528 ] = 8'h59;
  picture_data[ 2529 ] = 8'hE9;
  picture_data[ 2530 ] = 8'h49;
  picture_data[ 2531 ] = 8'hA9;
  picture_data[ 2532 ] = 8'h5A;
  picture_data[ 2533 ] = 8'h4C;
  picture_data[ 2534 ] = 8'h6A;
  picture_data[ 2535 ] = 8'hEE;
  picture_data[ 2536 ] = 8'h62;
  picture_data[ 2537 ] = 8'hCC;
  picture_data[ 2538 ] = 8'h4A;
  picture_data[ 2539 ] = 8'h29;
  picture_data[ 2540 ] = 8'h39;
  picture_data[ 2541 ] = 8'hC6;
  picture_data[ 2542 ] = 8'h62;
  picture_data[ 2543 ] = 8'hEB;
  picture_data[ 2544 ] = 8'h62;
  picture_data[ 2545 ] = 8'hCB;
  picture_data[ 2546 ] = 8'h5A;
  picture_data[ 2547 ] = 8'h69;
  picture_data[ 2548 ] = 8'h62;
  picture_data[ 2549 ] = 8'hA9;
  picture_data[ 2550 ] = 8'h41;
  picture_data[ 2551 ] = 8'hA5;
  picture_data[ 2552 ] = 8'h41;
  picture_data[ 2553 ] = 8'h83;
  picture_data[ 2554 ] = 8'h39;
  picture_data[ 2555 ] = 8'h42;
  picture_data[ 2556 ] = 8'h5A;
  picture_data[ 2557 ] = 8'h04;
  picture_data[ 2558 ] = 8'h72;
  picture_data[ 2559 ] = 8'h66;
  picture_data[ 2560 ] = 8'h8A;
  picture_data[ 2561 ] = 8'hA7;
  picture_data[ 2562 ] = 8'h82;
  picture_data[ 2563 ] = 8'h25;
  picture_data[ 2564 ] = 8'h81;
  picture_data[ 2565 ] = 8'hE5;
  picture_data[ 2566 ] = 8'h71;
  picture_data[ 2567 ] = 8'h63;
  picture_data[ 2568 ] = 8'hA3;
  picture_data[ 2569 ] = 8'hCB;
  picture_data[ 2570 ] = 8'hBD;
  picture_data[ 2571 ] = 8'h31;
  picture_data[ 2572 ] = 8'hB4;
  picture_data[ 2573 ] = 8'hCF;
  picture_data[ 2574 ] = 8'hB4;
  picture_data[ 2575 ] = 8'hEF;
  picture_data[ 2576 ] = 8'hB4;
  picture_data[ 2577 ] = 8'hEF;
  picture_data[ 2578 ] = 8'hBD;
  picture_data[ 2579 ] = 8'h31;
  picture_data[ 2580 ] = 8'hF7;
  picture_data[ 2581 ] = 8'h38;
  picture_data[ 2582 ] = 8'hDE;
  picture_data[ 2583 ] = 8'hD6;
  picture_data[ 2584 ] = 8'h19;
  picture_data[ 2585 ] = 8'h23;
  picture_data[ 2586 ] = 8'h08;
  picture_data[ 2587 ] = 8'hA1;
  picture_data[ 2588 ] = 8'h00;
  picture_data[ 2589 ] = 8'h81;
  picture_data[ 2590 ] = 8'h00;
  picture_data[ 2591 ] = 8'hA2;
  picture_data[ 2592 ] = 8'h00;
  picture_data[ 2593 ] = 8'h82;
  picture_data[ 2594 ] = 8'h08;
  picture_data[ 2595 ] = 8'hA2;
  picture_data[ 2596 ] = 8'h10;
  picture_data[ 2597 ] = 8'hE2;
  picture_data[ 2598 ] = 8'h19;
  picture_data[ 2599 ] = 8'h02;
  picture_data[ 2600 ] = 8'h18;
  picture_data[ 2601 ] = 8'hE2;
  picture_data[ 2602 ] = 8'h29;
  picture_data[ 2603 ] = 8'h85;
  picture_data[ 2604 ] = 8'h29;
  picture_data[ 2605 ] = 8'h65;
  picture_data[ 2606 ] = 8'h29;
  picture_data[ 2607 ] = 8'h24;
  picture_data[ 2608 ] = 8'h31;
  picture_data[ 2609 ] = 8'h23;
  picture_data[ 2610 ] = 8'h28;
  picture_data[ 2611 ] = 8'hA0;
  picture_data[ 2612 ] = 8'h9B;
  picture_data[ 2613 ] = 8'hC6;
  picture_data[ 2614 ] = 8'hF6;
  picture_data[ 2615 ] = 8'h4D;
  picture_data[ 2616 ] = 8'hCD;
  picture_data[ 2617 ] = 8'h07;
  picture_data[ 2618 ] = 8'hEE;
  picture_data[ 2619 ] = 8'h2E;
  picture_data[ 2620 ] = 8'h59;
  picture_data[ 2621 ] = 8'hA2;
  picture_data[ 2622 ] = 8'h20;
  picture_data[ 2623 ] = 8'h80;
  picture_data[ 2624 ] = 8'h29;
  picture_data[ 2625 ] = 8'h04;
  picture_data[ 2626 ] = 8'h10;
  picture_data[ 2627 ] = 8'h82;
  picture_data[ 2628 ] = 8'h10;
  picture_data[ 2629 ] = 8'hA2;
  picture_data[ 2630 ] = 8'h10;
  picture_data[ 2631 ] = 8'hC2;
  picture_data[ 2632 ] = 8'h10;
  picture_data[ 2633 ] = 8'hA0;
  picture_data[ 2634 ] = 8'h10;
  picture_data[ 2635 ] = 8'hE1;
  picture_data[ 2636 ] = 8'h21;
  picture_data[ 2637 ] = 8'h43;
  picture_data[ 2638 ] = 8'h19;
  picture_data[ 2639 ] = 8'h24;
  picture_data[ 2640 ] = 8'h29;
  picture_data[ 2641 ] = 8'hA8;
  picture_data[ 2642 ] = 8'h29;
  picture_data[ 2643 ] = 8'hC8;
  picture_data[ 2644 ] = 8'h19;
  picture_data[ 2645 ] = 8'h65;
  picture_data[ 2646 ] = 8'h32;
  picture_data[ 2647 ] = 8'h07;
  picture_data[ 2648 ] = 8'h31;
  picture_data[ 2649 ] = 8'hE8;
  picture_data[ 2650 ] = 8'h31;
  picture_data[ 2651 ] = 8'hC8;
  picture_data[ 2652 ] = 8'h21;
  picture_data[ 2653 ] = 8'h45;
  picture_data[ 2654 ] = 8'h21;
  picture_data[ 2655 ] = 8'h04;
  picture_data[ 2656 ] = 8'h18;
  picture_data[ 2657 ] = 8'hA2;
  picture_data[ 2658 ] = 8'h20;
  picture_data[ 2659 ] = 8'hA2;
  picture_data[ 2660 ] = 8'h28;
  picture_data[ 2661 ] = 8'hC3;
  picture_data[ 2662 ] = 8'h31;
  picture_data[ 2663 ] = 8'h04;
  picture_data[ 2664 ] = 8'h20;
  picture_data[ 2665 ] = 8'h82;
  picture_data[ 2666 ] = 8'h30;
  picture_data[ 2667 ] = 8'hC2;
  picture_data[ 2668 ] = 8'h41;
  picture_data[ 2669 ] = 8'h64;
  picture_data[ 2670 ] = 8'h6A;
  picture_data[ 2671 ] = 8'h88;
  picture_data[ 2672 ] = 8'h7B;
  picture_data[ 2673 ] = 8'h4B;
  picture_data[ 2674 ] = 8'h6A;
  picture_data[ 2675 ] = 8'hA9;
  picture_data[ 2676 ] = 8'h41;
  picture_data[ 2677 ] = 8'h85;
  picture_data[ 2678 ] = 8'h38;
  picture_data[ 2679 ] = 8'hE4;
  picture_data[ 2680 ] = 8'h49;
  picture_data[ 2681 ] = 8'h88;
  picture_data[ 2682 ] = 8'h72;
  picture_data[ 2683 ] = 8'hAD;
  picture_data[ 2684 ] = 8'h6A;
  picture_data[ 2685 ] = 8'hAD;
  picture_data[ 2686 ] = 8'h62;
  picture_data[ 2687 ] = 8'h8C;
  picture_data[ 2688 ] = 8'h62;
  picture_data[ 2689 ] = 8'hCC;
  picture_data[ 2690 ] = 8'h41;
  picture_data[ 2691 ] = 8'hE7;
  picture_data[ 2692 ] = 8'h42;
  picture_data[ 2693 ] = 8'h27;
  picture_data[ 2694 ] = 8'h4A;
  picture_data[ 2695 ] = 8'h48;
  picture_data[ 2696 ] = 8'h42;
  picture_data[ 2697 ] = 8'h08;
  picture_data[ 2698 ] = 8'h42;
  picture_data[ 2699 ] = 8'h08;
  picture_data[ 2700 ] = 8'h5A;
  picture_data[ 2701 ] = 8'h69;
  picture_data[ 2702 ] = 8'h5A;
  picture_data[ 2703 ] = 8'h68;
  picture_data[ 2704 ] = 8'h28;
  picture_data[ 2705 ] = 8'hC0;
  picture_data[ 2706 ] = 8'h59;
  picture_data[ 2707 ] = 8'hE4;
  picture_data[ 2708 ] = 8'h6A;
  picture_data[ 2709 ] = 8'h46;
  picture_data[ 2710 ] = 8'h6A;
  picture_data[ 2711 ] = 8'h05;
  picture_data[ 2712 ] = 8'h7A;
  picture_data[ 2713 ] = 8'h05;
  picture_data[ 2714 ] = 8'h79;
  picture_data[ 2715 ] = 8'h83;
  picture_data[ 2716 ] = 8'h89;
  picture_data[ 2717 ] = 8'hA4;
  picture_data[ 2718 ] = 8'h79;
  picture_data[ 2719 ] = 8'hA4;
  picture_data[ 2720 ] = 8'h93;
  picture_data[ 2721 ] = 8'h29;
  picture_data[ 2722 ] = 8'hBD;
  picture_data[ 2723 ] = 8'h10;
  picture_data[ 2724 ] = 8'hB5;
  picture_data[ 2725 ] = 8'h10;
  picture_data[ 2726 ] = 8'hB4;
  picture_data[ 2727 ] = 8'hF0;
  picture_data[ 2728 ] = 8'hB4;
  picture_data[ 2729 ] = 8'hF0;
  picture_data[ 2730 ] = 8'hBD;
  picture_data[ 2731 ] = 8'h30;
  picture_data[ 2732 ] = 8'hEF;
  picture_data[ 2733 ] = 8'h17;
  picture_data[ 2734 ] = 8'hDE;
  picture_data[ 2735 ] = 8'hD6;
  picture_data[ 2736 ] = 8'h08;
  picture_data[ 2737 ] = 8'hC2;
  picture_data[ 2738 ] = 8'h08;
  picture_data[ 2739 ] = 8'hA1;
  picture_data[ 2740 ] = 8'h00;
  picture_data[ 2741 ] = 8'hA1;
  picture_data[ 2742 ] = 8'h08;
  picture_data[ 2743 ] = 8'hE2;
  picture_data[ 2744 ] = 8'h19;
  picture_data[ 2745 ] = 8'h24;
  picture_data[ 2746 ] = 8'h10;
  picture_data[ 2747 ] = 8'hE3;
  picture_data[ 2748 ] = 8'h10;
  picture_data[ 2749 ] = 8'hC1;
  picture_data[ 2750 ] = 8'h19;
  picture_data[ 2751 ] = 8'h02;
  picture_data[ 2752 ] = 8'h21;
  picture_data[ 2753 ] = 8'h43;
  picture_data[ 2754 ] = 8'h29;
  picture_data[ 2755 ] = 8'h64;
  picture_data[ 2756 ] = 8'h18;
  picture_data[ 2757 ] = 8'hE3;
  picture_data[ 2758 ] = 8'h20;
  picture_data[ 2759 ] = 8'hE4;
  picture_data[ 2760 ] = 8'h28;
  picture_data[ 2761 ] = 8'hE3;
  picture_data[ 2762 ] = 8'h28;
  picture_data[ 2763 ] = 8'hA0;
  picture_data[ 2764 ] = 8'h41;
  picture_data[ 2765 ] = 8'h40;
  picture_data[ 2766 ] = 8'hC5;
  picture_data[ 2767 ] = 8'h0B;
  picture_data[ 2768 ] = 8'hE5;
  picture_data[ 2769 ] = 8'hEE;
  picture_data[ 2770 ] = 8'h8B;
  picture_data[ 2771 ] = 8'h45;
  picture_data[ 2772 ] = 8'h30;
  picture_data[ 2773 ] = 8'hC0;
  picture_data[ 2774 ] = 8'h28;
  picture_data[ 2775 ] = 8'hC1;
  picture_data[ 2776 ] = 8'h20;
  picture_data[ 2777 ] = 8'hE2;
  picture_data[ 2778 ] = 8'h31;
  picture_data[ 2779 ] = 8'h85;
  picture_data[ 2780 ] = 8'h18;
  picture_data[ 2781 ] = 8'hA1;
  picture_data[ 2782 ] = 8'h21;
  picture_data[ 2783 ] = 8'h02;
  picture_data[ 2784 ] = 8'h31;
  picture_data[ 2785 ] = 8'hA4;
  picture_data[ 2786 ] = 8'h39;
  picture_data[ 2787 ] = 8'hC4;
  picture_data[ 2788 ] = 8'h31;
  picture_data[ 2789 ] = 8'h84;
  picture_data[ 2790 ] = 8'h29;
  picture_data[ 2791 ] = 8'h85;
  picture_data[ 2792 ] = 8'h31;
  picture_data[ 2793 ] = 8'hA8;
  picture_data[ 2794 ] = 8'h29;
  picture_data[ 2795 ] = 8'h88;
  picture_data[ 2796 ] = 8'h19;
  picture_data[ 2797 ] = 8'h46;
  picture_data[ 2798 ] = 8'h29;
  picture_data[ 2799 ] = 8'hA7;
  picture_data[ 2800 ] = 8'h29;
  picture_data[ 2801 ] = 8'hA8;
  picture_data[ 2802 ] = 8'h31;
  picture_data[ 2803 ] = 8'hC9;
  picture_data[ 2804 ] = 8'h18;
  picture_data[ 2805 ] = 8'hC4;
  picture_data[ 2806 ] = 8'h10;
  picture_data[ 2807 ] = 8'h63;
  picture_data[ 2808 ] = 8'h18;
  picture_data[ 2809 ] = 8'h83;
  picture_data[ 2810 ] = 8'h18;
  picture_data[ 2811 ] = 8'h83;
  picture_data[ 2812 ] = 8'h20;
  picture_data[ 2813 ] = 8'hA4;
  picture_data[ 2814 ] = 8'h30;
  picture_data[ 2815 ] = 8'hE5;
  picture_data[ 2816 ] = 8'h30;
  picture_data[ 2817 ] = 8'hE5;
  picture_data[ 2818 ] = 8'h20;
  picture_data[ 2819 ] = 8'h42;
  picture_data[ 2820 ] = 8'h28;
  picture_data[ 2821 ] = 8'h82;
  picture_data[ 2822 ] = 8'h28;
  picture_data[ 2823 ] = 8'h82;
  picture_data[ 2824 ] = 8'h30;
  picture_data[ 2825 ] = 8'hC2;
  picture_data[ 2826 ] = 8'h28;
  picture_data[ 2827 ] = 8'h82;
  picture_data[ 2828 ] = 8'h20;
  picture_data[ 2829 ] = 8'h41;
  picture_data[ 2830 ] = 8'h41;
  picture_data[ 2831 ] = 8'h66;
  picture_data[ 2832 ] = 8'h62;
  picture_data[ 2833 ] = 8'h4B;
  picture_data[ 2834 ] = 8'h62;
  picture_data[ 2835 ] = 8'h6C;
  picture_data[ 2836 ] = 8'h72;
  picture_data[ 2837 ] = 8'hEE;
  picture_data[ 2838 ] = 8'h62;
  picture_data[ 2839 ] = 8'h8C;
  picture_data[ 2840 ] = 8'h41;
  picture_data[ 2841 ] = 8'hE7;
  picture_data[ 2842 ] = 8'h42;
  picture_data[ 2843 ] = 8'h07;
  picture_data[ 2844 ] = 8'h39;
  picture_data[ 2845 ] = 8'hC6;
  picture_data[ 2846 ] = 8'h39;
  picture_data[ 2847 ] = 8'hE6;
  picture_data[ 2848 ] = 8'h31;
  picture_data[ 2849 ] = 8'h85;
  picture_data[ 2850 ] = 8'h52;
  picture_data[ 2851 ] = 8'h8A;
  picture_data[ 2852 ] = 8'h52;
  picture_data[ 2853 ] = 8'h49;
  picture_data[ 2854 ] = 8'h52;
  picture_data[ 2855 ] = 8'h27;
  picture_data[ 2856 ] = 8'h39;
  picture_data[ 2857 ] = 8'h42;
  picture_data[ 2858 ] = 8'h5A;
  picture_data[ 2859 ] = 8'h25;
  picture_data[ 2860 ] = 8'h51;
  picture_data[ 2861 ] = 8'hC4;
  picture_data[ 2862 ] = 8'h51;
  picture_data[ 2863 ] = 8'h83;
  picture_data[ 2864 ] = 8'h61;
  picture_data[ 2865 ] = 8'hA4;
  picture_data[ 2866 ] = 8'h79;
  picture_data[ 2867 ] = 8'hC4;
  picture_data[ 2868 ] = 8'h79;
  picture_data[ 2869 ] = 8'hA4;
  picture_data[ 2870 ] = 8'h69;
  picture_data[ 2871 ] = 8'h63;
  picture_data[ 2872 ] = 8'h7A;
  picture_data[ 2873 ] = 8'hA7;
  picture_data[ 2874 ] = 8'hC5;
  picture_data[ 2875 ] = 8'h51;
  picture_data[ 2876 ] = 8'hAC;
  picture_data[ 2877 ] = 8'hCF;
  picture_data[ 2878 ] = 8'hB4;
  picture_data[ 2879 ] = 8'hEF;
  picture_data[ 2880 ] = 8'hB4;
  picture_data[ 2881 ] = 8'hEF;
  picture_data[ 2882 ] = 8'hB4;
  picture_data[ 2883 ] = 8'hEF;
  picture_data[ 2884 ] = 8'hEE;
  picture_data[ 2885 ] = 8'hD6;
  picture_data[ 2886 ] = 8'hF7;
  picture_data[ 2887 ] = 8'h17;
  picture_data[ 2888 ] = 8'h19;
  picture_data[ 2889 ] = 8'h23;
  picture_data[ 2890 ] = 8'h08;
  picture_data[ 2891 ] = 8'hC2;
  picture_data[ 2892 ] = 8'h08;
  picture_data[ 2893 ] = 8'hE2;
  picture_data[ 2894 ] = 8'h08;
  picture_data[ 2895 ] = 8'hE2;
  picture_data[ 2896 ] = 8'h00;
  picture_data[ 2897 ] = 8'hA1;
  picture_data[ 2898 ] = 8'h08;
  picture_data[ 2899 ] = 8'hA1;
  picture_data[ 2900 ] = 8'h08;
  picture_data[ 2901 ] = 8'hC1;
  picture_data[ 2902 ] = 8'h08;
  picture_data[ 2903 ] = 8'hA1;
  picture_data[ 2904 ] = 8'h10;
  picture_data[ 2905 ] = 8'hE2;
  picture_data[ 2906 ] = 8'h21;
  picture_data[ 2907 ] = 8'h64;
  picture_data[ 2908 ] = 8'h19;
  picture_data[ 2909 ] = 8'h44;
  picture_data[ 2910 ] = 8'h10;
  picture_data[ 2911 ] = 8'hC3;
  picture_data[ 2912 ] = 8'h10;
  picture_data[ 2913 ] = 8'h41;
  picture_data[ 2914 ] = 8'h18;
  picture_data[ 2915 ] = 8'h80;
  picture_data[ 2916 ] = 8'h31;
  picture_data[ 2917 ] = 8'h00;
  picture_data[ 2918 ] = 8'h30;
  picture_data[ 2919 ] = 8'hA0;
  picture_data[ 2920 ] = 8'h49;
  picture_data[ 2921 ] = 8'h60;
  picture_data[ 2922 ] = 8'h39;
  picture_data[ 2923 ] = 8'h00;
  picture_data[ 2924 ] = 8'h30;
  picture_data[ 2925 ] = 8'hC0;
  picture_data[ 2926 ] = 8'h20;
  picture_data[ 2927 ] = 8'h80;
  picture_data[ 2928 ] = 8'h31;
  picture_data[ 2929 ] = 8'h02;
  picture_data[ 2930 ] = 8'h5A;
  picture_data[ 2931 ] = 8'h88;
  picture_data[ 2932 ] = 8'h41;
  picture_data[ 2933 ] = 8'hA5;
  picture_data[ 2934 ] = 8'h62;
  picture_data[ 2935 ] = 8'hC9;
  picture_data[ 2936 ] = 8'h83;
  picture_data[ 2937 ] = 8'hCD;
  picture_data[ 2938 ] = 8'h73;
  picture_data[ 2939 ] = 8'h6B;
  picture_data[ 2940 ] = 8'h62;
  picture_data[ 2941 ] = 8'hE9;
  picture_data[ 2942 ] = 8'h62;
  picture_data[ 2943 ] = 8'hEA;
  picture_data[ 2944 ] = 8'h41;
  picture_data[ 2945 ] = 8'hEA;
  picture_data[ 2946 ] = 8'h31;
  picture_data[ 2947 ] = 8'hA9;
  picture_data[ 2948 ] = 8'h19;
  picture_data[ 2949 ] = 8'h25;
  picture_data[ 2950 ] = 8'h29;
  picture_data[ 2951 ] = 8'h87;
  picture_data[ 2952 ] = 8'h31;
  picture_data[ 2953 ] = 8'hA9;
  picture_data[ 2954 ] = 8'h29;
  picture_data[ 2955 ] = 8'h68;
  picture_data[ 2956 ] = 8'h21;
  picture_data[ 2957 ] = 8'h06;
  picture_data[ 2958 ] = 8'h20;
  picture_data[ 2959 ] = 8'hE5;
  picture_data[ 2960 ] = 8'h20;
  picture_data[ 2961 ] = 8'hC4;
  picture_data[ 2962 ] = 8'h20;
  picture_data[ 2963 ] = 8'hC5;
  picture_data[ 2964 ] = 8'h31;
  picture_data[ 2965 ] = 8'h06;
  picture_data[ 2966 ] = 8'h31;
  picture_data[ 2967 ] = 8'h27;
  picture_data[ 2968 ] = 8'h41;
  picture_data[ 2969 ] = 8'h68;
  picture_data[ 2970 ] = 8'h28;
  picture_data[ 2971 ] = 8'hA4;
  picture_data[ 2972 ] = 8'h30;
  picture_data[ 2973 ] = 8'hE4;
  picture_data[ 2974 ] = 8'h30;
  picture_data[ 2975 ] = 8'hC4;
  picture_data[ 2976 ] = 8'h39;
  picture_data[ 2977 ] = 8'h04;
  picture_data[ 2978 ] = 8'h38;
  picture_data[ 2979 ] = 8'hE4;
  picture_data[ 2980 ] = 8'h39;
  picture_data[ 2981 ] = 8'h05;
  picture_data[ 2982 ] = 8'h49;
  picture_data[ 2983 ] = 8'h87;
  picture_data[ 2984 ] = 8'h62;
  picture_data[ 2985 ] = 8'h6B;
  picture_data[ 2986 ] = 8'h62;
  picture_data[ 2987 ] = 8'h8B;
  picture_data[ 2988 ] = 8'h5A;
  picture_data[ 2989 ] = 8'h4A;
  picture_data[ 2990 ] = 8'h73;
  picture_data[ 2991 ] = 8'h4E;
  picture_data[ 2992 ] = 8'h52;
  picture_data[ 2993 ] = 8'h48;
  picture_data[ 2994 ] = 8'h29;
  picture_data[ 2995 ] = 8'h43;
  picture_data[ 2996 ] = 8'h39;
  picture_data[ 2997 ] = 8'hE6;
  picture_data[ 2998 ] = 8'h29;
  picture_data[ 2999 ] = 8'h64;
  picture_data[ 3000 ] = 8'h31;
  picture_data[ 3001 ] = 8'h85;
  picture_data[ 3002 ] = 8'h39;
  picture_data[ 3003 ] = 8'hC7;
  picture_data[ 3004 ] = 8'h29;
  picture_data[ 3005 ] = 8'h03;
  picture_data[ 3006 ] = 8'h41;
  picture_data[ 3007 ] = 8'h85;
  picture_data[ 3008 ] = 8'h49;
  picture_data[ 3009 ] = 8'hC4;
  picture_data[ 3010 ] = 8'h49;
  picture_data[ 3011 ] = 8'hC4;
  picture_data[ 3012 ] = 8'h5A;
  picture_data[ 3013 ] = 8'h05;
  picture_data[ 3014 ] = 8'h59;
  picture_data[ 3015 ] = 8'hC4;
  picture_data[ 3016 ] = 8'h6A;
  picture_data[ 3017 ] = 8'h04;
  picture_data[ 3018 ] = 8'h72;
  picture_data[ 3019 ] = 8'h04;
  picture_data[ 3020 ] = 8'h82;
  picture_data[ 3021 ] = 8'h25;
  picture_data[ 3022 ] = 8'h71;
  picture_data[ 3023 ] = 8'hA4;
  picture_data[ 3024 ] = 8'h61;
  picture_data[ 3025 ] = 8'hC3;
  picture_data[ 3026 ] = 8'hC5;
  picture_data[ 3027 ] = 8'h51;
  picture_data[ 3028 ] = 8'hB4;
  picture_data[ 3029 ] = 8'hEF;
  picture_data[ 3030 ] = 8'hAC;
  picture_data[ 3031 ] = 8'hEF;
  picture_data[ 3032 ] = 8'hB5;
  picture_data[ 3033 ] = 8'h0F;
  picture_data[ 3034 ] = 8'hB4;
  picture_data[ 3035 ] = 8'hEF;
  picture_data[ 3036 ] = 8'hE6;
  picture_data[ 3037 ] = 8'h95;
  picture_data[ 3038 ] = 8'hF7;
  picture_data[ 3039 ] = 8'h17;
  picture_data[ 3040 ] = 8'h19;
  picture_data[ 3041 ] = 8'h23;
  picture_data[ 3042 ] = 8'h19;
  picture_data[ 3043 ] = 8'h44;
  picture_data[ 3044 ] = 8'h08;
  picture_data[ 3045 ] = 8'hE2;
  picture_data[ 3046 ] = 8'h00;
  picture_data[ 3047 ] = 8'h81;
  picture_data[ 3048 ] = 8'h00;
  picture_data[ 3049 ] = 8'h81;
  picture_data[ 3050 ] = 8'h00;
  picture_data[ 3051 ] = 8'h81;
  picture_data[ 3052 ] = 8'h00;
  picture_data[ 3053 ] = 8'h80;
  picture_data[ 3054 ] = 8'h10;
  picture_data[ 3055 ] = 8'hE1;
  picture_data[ 3056 ] = 8'h08;
  picture_data[ 3057 ] = 8'hA1;
  picture_data[ 3058 ] = 8'h08;
  picture_data[ 3059 ] = 8'hC2;
  picture_data[ 3060 ] = 8'h19;
  picture_data[ 3061 ] = 8'h24;
  picture_data[ 3062 ] = 8'h08;
  picture_data[ 3063 ] = 8'hC2;
  picture_data[ 3064 ] = 8'h19;
  picture_data[ 3065 ] = 8'h04;
  picture_data[ 3066 ] = 8'h29;
  picture_data[ 3067 ] = 8'h44;
  picture_data[ 3068 ] = 8'h31;
  picture_data[ 3069 ] = 8'h21;
  picture_data[ 3070 ] = 8'h28;
  picture_data[ 3071 ] = 8'hC0;
  picture_data[ 3072 ] = 8'h28;
  picture_data[ 3073 ] = 8'hC0;
  picture_data[ 3074 ] = 8'h31;
  picture_data[ 3075 ] = 8'h01;
  picture_data[ 3076 ] = 8'h41;
  picture_data[ 3077 ] = 8'h83;
  picture_data[ 3078 ] = 8'h5A;
  picture_data[ 3079 ] = 8'h26;
  picture_data[ 3080 ] = 8'h6A;
  picture_data[ 3081 ] = 8'hA8;
  picture_data[ 3082 ] = 8'h83;
  picture_data[ 3083 ] = 8'h8B;
  picture_data[ 3084 ] = 8'h7B;
  picture_data[ 3085 ] = 8'h2B;
  picture_data[ 3086 ] = 8'h83;
  picture_data[ 3087 ] = 8'h8C;
  picture_data[ 3088 ] = 8'h83;
  picture_data[ 3089 ] = 8'h6C;
  picture_data[ 3090 ] = 8'h62;
  picture_data[ 3091 ] = 8'h67;
  picture_data[ 3092 ] = 8'h73;
  picture_data[ 3093 ] = 8'h2A;
  picture_data[ 3094 ] = 8'h73;
  picture_data[ 3095 ] = 8'h0B;
  picture_data[ 3096 ] = 8'h39;
  picture_data[ 3097 ] = 8'h87;
  picture_data[ 3098 ] = 8'h39;
  picture_data[ 3099 ] = 8'h88;
  picture_data[ 3100 ] = 8'h10;
  picture_data[ 3101 ] = 8'hA3;
  picture_data[ 3102 ] = 8'h31;
  picture_data[ 3103 ] = 8'h87;
  picture_data[ 3104 ] = 8'h31;
  picture_data[ 3105 ] = 8'h67;
  picture_data[ 3106 ] = 8'h29;
  picture_data[ 3107 ] = 8'h47;
  picture_data[ 3108 ] = 8'h21;
  picture_data[ 3109 ] = 8'h05;
  picture_data[ 3110 ] = 8'h18;
  picture_data[ 3111 ] = 8'hA4;
  picture_data[ 3112 ] = 8'h20;
  picture_data[ 3113 ] = 8'hE5;
  picture_data[ 3114 ] = 8'h20;
  picture_data[ 3115 ] = 8'hA4;
  picture_data[ 3116 ] = 8'h18;
  picture_data[ 3117 ] = 8'h63;
  picture_data[ 3118 ] = 8'h39;
  picture_data[ 3119 ] = 8'h68;
  picture_data[ 3120 ] = 8'h39;
  picture_data[ 3121 ] = 8'h27;
  picture_data[ 3122 ] = 8'h51;
  picture_data[ 3123 ] = 8'hC9;
  picture_data[ 3124 ] = 8'h30;
  picture_data[ 3125 ] = 8'hE4;
  picture_data[ 3126 ] = 8'h30;
  picture_data[ 3127 ] = 8'hE4;
  picture_data[ 3128 ] = 8'h49;
  picture_data[ 3129 ] = 8'h86;
  picture_data[ 3130 ] = 8'h51;
  picture_data[ 3131 ] = 8'hE8;
  picture_data[ 3132 ] = 8'h49;
  picture_data[ 3133 ] = 8'hA7;
  picture_data[ 3134 ] = 8'h41;
  picture_data[ 3135 ] = 8'h66;
  picture_data[ 3136 ] = 8'h52;
  picture_data[ 3137 ] = 8'h09;
  picture_data[ 3138 ] = 8'h5A;
  picture_data[ 3139 ] = 8'h4A;
  picture_data[ 3140 ] = 8'h5A;
  picture_data[ 3141 ] = 8'h8A;
  picture_data[ 3142 ] = 8'h52;
  picture_data[ 3143 ] = 8'h28;
  picture_data[ 3144 ] = 8'h5A;
  picture_data[ 3145 ] = 8'hCA;
  picture_data[ 3146 ] = 8'h29;
  picture_data[ 3147 ] = 8'h64;
  picture_data[ 3148 ] = 8'h29;
  picture_data[ 3149 ] = 8'h64;
  picture_data[ 3150 ] = 8'h31;
  picture_data[ 3151 ] = 8'h84;
  picture_data[ 3152 ] = 8'h42;
  picture_data[ 3153 ] = 8'h07;
  picture_data[ 3154 ] = 8'h39;
  picture_data[ 3155 ] = 8'hC6;
  picture_data[ 3156 ] = 8'h4A;
  picture_data[ 3157 ] = 8'h27;
  picture_data[ 3158 ] = 8'h52;
  picture_data[ 3159 ] = 8'h27;
  picture_data[ 3160 ] = 8'h52;
  picture_data[ 3161 ] = 8'h26;
  picture_data[ 3162 ] = 8'h73;
  picture_data[ 3163 ] = 8'h29;
  picture_data[ 3164 ] = 8'h49;
  picture_data[ 3165 ] = 8'hC4;
  picture_data[ 3166 ] = 8'h49;
  picture_data[ 3167 ] = 8'hA3;
  picture_data[ 3168 ] = 8'h6A;
  picture_data[ 3169 ] = 8'h24;
  picture_data[ 3170 ] = 8'h72;
  picture_data[ 3171 ] = 8'h03;
  picture_data[ 3172 ] = 8'h69;
  picture_data[ 3173 ] = 8'h62;
  picture_data[ 3174 ] = 8'h79;
  picture_data[ 3175 ] = 8'hE4;
  picture_data[ 3176 ] = 8'h61;
  picture_data[ 3177 ] = 8'hA2;
  picture_data[ 3178 ] = 8'hBC;
  picture_data[ 3179 ] = 8'hCE;
  picture_data[ 3180 ] = 8'hB5;
  picture_data[ 3181 ] = 8'h0F;
  picture_data[ 3182 ] = 8'hB5;
  picture_data[ 3183 ] = 8'h50;
  picture_data[ 3184 ] = 8'hAD;
  picture_data[ 3185 ] = 8'h2F;
  picture_data[ 3186 ] = 8'hAC;
  picture_data[ 3187 ] = 8'hEF;
  picture_data[ 3188 ] = 8'hD6;
  picture_data[ 3189 ] = 8'h34;
  picture_data[ 3190 ] = 8'hF7;
  picture_data[ 3191 ] = 8'h18;
  picture_data[ 3192 ] = 8'h08;
  picture_data[ 3193 ] = 8'hC2;
  picture_data[ 3194 ] = 8'h00;
  picture_data[ 3195 ] = 8'hA2;
  picture_data[ 3196 ] = 8'h08;
  picture_data[ 3197 ] = 8'hE2;
  picture_data[ 3198 ] = 8'h11;
  picture_data[ 3199 ] = 8'h03;
  picture_data[ 3200 ] = 8'h08;
  picture_data[ 3201 ] = 8'hA2;
  picture_data[ 3202 ] = 8'h00;
  picture_data[ 3203 ] = 8'hA1;
  picture_data[ 3204 ] = 8'h08;
  picture_data[ 3205 ] = 8'hC2;
  picture_data[ 3206 ] = 8'h10;
  picture_data[ 3207 ] = 8'hC2;
  picture_data[ 3208 ] = 8'h11;
  picture_data[ 3209 ] = 8'h02;
  picture_data[ 3210 ] = 8'h11;
  picture_data[ 3211 ] = 8'h23;
  picture_data[ 3212 ] = 8'h11;
  picture_data[ 3213 ] = 8'h02;
  picture_data[ 3214 ] = 8'h21;
  picture_data[ 3215 ] = 8'h64;
  picture_data[ 3216 ] = 8'h29;
  picture_data[ 3217 ] = 8'h65;
  picture_data[ 3218 ] = 8'h29;
  picture_data[ 3219 ] = 8'h64;
  picture_data[ 3220 ] = 8'h39;
  picture_data[ 3221 ] = 8'h84;
  picture_data[ 3222 ] = 8'h29;
  picture_data[ 3223 ] = 8'h02;
  picture_data[ 3224 ] = 8'h31;
  picture_data[ 3225 ] = 8'h22;
  picture_data[ 3226 ] = 8'h39;
  picture_data[ 3227 ] = 8'h43;
  picture_data[ 3228 ] = 8'h62;
  picture_data[ 3229 ] = 8'h68;
  picture_data[ 3230 ] = 8'h7B;
  picture_data[ 3231 ] = 8'h2A;
  picture_data[ 3232 ] = 8'h83;
  picture_data[ 3233 ] = 8'h6A;
  picture_data[ 3234 ] = 8'h8B;
  picture_data[ 3235 ] = 8'h8B;
  picture_data[ 3236 ] = 8'h83;
  picture_data[ 3237 ] = 8'h2A;
  picture_data[ 3238 ] = 8'h7B;
  picture_data[ 3239 ] = 8'h2B;
  picture_data[ 3240 ] = 8'h72;
  picture_data[ 3241 ] = 8'hC9;
  picture_data[ 3242 ] = 8'h51;
  picture_data[ 3243 ] = 8'hE6;
  picture_data[ 3244 ] = 8'h6A;
  picture_data[ 3245 ] = 8'hA9;
  picture_data[ 3246 ] = 8'h72;
  picture_data[ 3247 ] = 8'hEA;
  picture_data[ 3248 ] = 8'h41;
  picture_data[ 3249 ] = 8'h87;
  picture_data[ 3250 ] = 8'h31;
  picture_data[ 3251 ] = 8'h67;
  picture_data[ 3252 ] = 8'h20;
  picture_data[ 3253 ] = 8'hE4;
  picture_data[ 3254 ] = 8'h31;
  picture_data[ 3255 ] = 8'h66;
  picture_data[ 3256 ] = 8'h31;
  picture_data[ 3257 ] = 8'h87;
  picture_data[ 3258 ] = 8'h20;
  picture_data[ 3259 ] = 8'hC4;
  picture_data[ 3260 ] = 8'h20;
  picture_data[ 3261 ] = 8'hE4;
  picture_data[ 3262 ] = 8'h20;
  picture_data[ 3263 ] = 8'hE4;
  picture_data[ 3264 ] = 8'h31;
  picture_data[ 3265 ] = 8'h25;
  picture_data[ 3266 ] = 8'h31;
  picture_data[ 3267 ] = 8'h25;
  picture_data[ 3268 ] = 8'h28;
  picture_data[ 3269 ] = 8'hE5;
  picture_data[ 3270 ] = 8'h39;
  picture_data[ 3271 ] = 8'h88;
  picture_data[ 3272 ] = 8'h20;
  picture_data[ 3273 ] = 8'h84;
  picture_data[ 3274 ] = 8'h49;
  picture_data[ 3275 ] = 8'hC8;
  picture_data[ 3276 ] = 8'h49;
  picture_data[ 3277 ] = 8'hA7;
  picture_data[ 3278 ] = 8'h30;
  picture_data[ 3279 ] = 8'hE3;
  picture_data[ 3280 ] = 8'h41;
  picture_data[ 3281 ] = 8'h65;
  picture_data[ 3282 ] = 8'h51;
  picture_data[ 3283 ] = 8'hE7;
  picture_data[ 3284 ] = 8'h41;
  picture_data[ 3285 ] = 8'h65;
  picture_data[ 3286 ] = 8'h49;
  picture_data[ 3287 ] = 8'hA6;
  picture_data[ 3288 ] = 8'h49;
  picture_data[ 3289 ] = 8'hE7;
  picture_data[ 3290 ] = 8'h4A;
  picture_data[ 3291 ] = 8'h08;
  picture_data[ 3292 ] = 8'h41;
  picture_data[ 3293 ] = 8'hC7;
  picture_data[ 3294 ] = 8'h29;
  picture_data[ 3295 ] = 8'h03;
  picture_data[ 3296 ] = 8'h52;
  picture_data[ 3297 ] = 8'h68;
  picture_data[ 3298 ] = 8'h39;
  picture_data[ 3299 ] = 8'hA4;
  picture_data[ 3300 ] = 8'h29;
  picture_data[ 3301 ] = 8'h63;
  picture_data[ 3302 ] = 8'h29;
  picture_data[ 3303 ] = 8'h84;
  picture_data[ 3304 ] = 8'h31;
  picture_data[ 3305 ] = 8'hA5;
  picture_data[ 3306 ] = 8'h41;
  picture_data[ 3307 ] = 8'hE6;
  picture_data[ 3308 ] = 8'h52;
  picture_data[ 3309 ] = 8'h89;
  picture_data[ 3310 ] = 8'h5A;
  picture_data[ 3311 ] = 8'h88;
  picture_data[ 3312 ] = 8'h39;
  picture_data[ 3313 ] = 8'hA4;
  picture_data[ 3314 ] = 8'h62;
  picture_data[ 3315 ] = 8'hE8;
  picture_data[ 3316 ] = 8'h6B;
  picture_data[ 3317 ] = 8'h09;
  picture_data[ 3318 ] = 8'h5A;
  picture_data[ 3319 ] = 8'h25;
  picture_data[ 3320 ] = 8'h62;
  picture_data[ 3321 ] = 8'h24;
  picture_data[ 3322 ] = 8'h72;
  picture_data[ 3323 ] = 8'h23;
  picture_data[ 3324 ] = 8'h72;
  picture_data[ 3325 ] = 8'h03;
  picture_data[ 3326 ] = 8'h82;
  picture_data[ 3327 ] = 8'h65;
  picture_data[ 3328 ] = 8'h9B;
  picture_data[ 3329 ] = 8'h48;
  picture_data[ 3330 ] = 8'h8B;
  picture_data[ 3331 ] = 8'h28;
  picture_data[ 3332 ] = 8'hB4;
  picture_data[ 3333 ] = 8'hEE;
  picture_data[ 3334 ] = 8'hAC;
  picture_data[ 3335 ] = 8'hEE;
  picture_data[ 3336 ] = 8'hAD;
  picture_data[ 3337 ] = 8'h0F;
  picture_data[ 3338 ] = 8'hAD;
  picture_data[ 3339 ] = 8'h2F;
  picture_data[ 3340 ] = 8'hD6;
  picture_data[ 3341 ] = 8'h55;
  picture_data[ 3342 ] = 8'hFF;
  picture_data[ 3343 ] = 8'h9A;
  picture_data[ 3344 ] = 8'h08;
  picture_data[ 3345 ] = 8'hA2;
  picture_data[ 3346 ] = 8'h08;
  picture_data[ 3347 ] = 8'hA2;
  picture_data[ 3348 ] = 8'h00;
  picture_data[ 3349 ] = 8'hA2;
  picture_data[ 3350 ] = 8'h08;
  picture_data[ 3351 ] = 8'hE3;
  picture_data[ 3352 ] = 8'h08;
  picture_data[ 3353 ] = 8'hE3;
  picture_data[ 3354 ] = 8'h00;
  picture_data[ 3355 ] = 8'h82;
  picture_data[ 3356 ] = 8'h00;
  picture_data[ 3357 ] = 8'h61;
  picture_data[ 3358 ] = 8'h08;
  picture_data[ 3359 ] = 8'hC2;
  picture_data[ 3360 ] = 8'h08;
  picture_data[ 3361 ] = 8'hC2;
  picture_data[ 3362 ] = 8'h10;
  picture_data[ 3363 ] = 8'hE2;
  picture_data[ 3364 ] = 8'h11;
  picture_data[ 3365 ] = 8'h02;
  picture_data[ 3366 ] = 8'h21;
  picture_data[ 3367 ] = 8'hA4;
  picture_data[ 3368 ] = 8'h3A;
  picture_data[ 3369 ] = 8'h47;
  picture_data[ 3370 ] = 8'h21;
  picture_data[ 3371 ] = 8'h23;
  picture_data[ 3372 ] = 8'h39;
  picture_data[ 3373 ] = 8'hE6;
  picture_data[ 3374 ] = 8'h39;
  picture_data[ 3375 ] = 8'h84;
  picture_data[ 3376 ] = 8'h52;
  picture_data[ 3377 ] = 8'h67;
  picture_data[ 3378 ] = 8'h52;
  picture_data[ 3379 ] = 8'h47;
  picture_data[ 3380 ] = 8'h72;
  picture_data[ 3381 ] = 8'hEA;
  picture_data[ 3382 ] = 8'h8B;
  picture_data[ 3383 ] = 8'h8C;
  picture_data[ 3384 ] = 8'h7B;
  picture_data[ 3385 ] = 8'h09;
  picture_data[ 3386 ] = 8'h72;
  picture_data[ 3387 ] = 8'hA7;
  picture_data[ 3388 ] = 8'h83;
  picture_data[ 3389 ] = 8'h2A;
  picture_data[ 3390 ] = 8'h8B;
  picture_data[ 3391 ] = 8'h6C;
  picture_data[ 3392 ] = 8'h7B;
  picture_data[ 3393 ] = 8'h0B;
  picture_data[ 3394 ] = 8'h62;
  picture_data[ 3395 ] = 8'h48;
  picture_data[ 3396 ] = 8'h6A;
  picture_data[ 3397 ] = 8'hA9;
  picture_data[ 3398 ] = 8'h7B;
  picture_data[ 3399 ] = 8'h0B;
  picture_data[ 3400 ] = 8'h62;
  picture_data[ 3401 ] = 8'h69;
  picture_data[ 3402 ] = 8'h28;
  picture_data[ 3403 ] = 8'hE4;
  picture_data[ 3404 ] = 8'h29;
  picture_data[ 3405 ] = 8'h24;
  picture_data[ 3406 ] = 8'h29;
  picture_data[ 3407 ] = 8'h24;
  picture_data[ 3408 ] = 8'h29;
  picture_data[ 3409 ] = 8'h04;
  picture_data[ 3410 ] = 8'h29;
  picture_data[ 3411 ] = 8'h04;
  picture_data[ 3412 ] = 8'h28;
  picture_data[ 3413 ] = 8'hE4;
  picture_data[ 3414 ] = 8'h20;
  picture_data[ 3415 ] = 8'hE3;
  picture_data[ 3416 ] = 8'h41;
  picture_data[ 3417 ] = 8'hC7;
  picture_data[ 3418 ] = 8'h39;
  picture_data[ 3419 ] = 8'hA7;
  picture_data[ 3420 ] = 8'h29;
  picture_data[ 3421 ] = 8'h05;
  picture_data[ 3422 ] = 8'h39;
  picture_data[ 3423 ] = 8'h87;
  picture_data[ 3424 ] = 8'h39;
  picture_data[ 3425 ] = 8'h67;
  picture_data[ 3426 ] = 8'h41;
  picture_data[ 3427 ] = 8'hA7;
  picture_data[ 3428 ] = 8'h49;
  picture_data[ 3429 ] = 8'hC7;
  picture_data[ 3430 ] = 8'h39;
  picture_data[ 3431 ] = 8'h65;
  picture_data[ 3432 ] = 8'h49;
  picture_data[ 3433 ] = 8'hA5;
  picture_data[ 3434 ] = 8'h49;
  picture_data[ 3435 ] = 8'hC6;
  picture_data[ 3436 ] = 8'h41;
  picture_data[ 3437 ] = 8'h85;
  picture_data[ 3438 ] = 8'h52;
  picture_data[ 3439 ] = 8'h07;
  picture_data[ 3440 ] = 8'h4A;
  picture_data[ 3441 ] = 8'h07;
  picture_data[ 3442 ] = 8'h39;
  picture_data[ 3443 ] = 8'hA5;
  picture_data[ 3444 ] = 8'h31;
  picture_data[ 3445 ] = 8'h64;
  picture_data[ 3446 ] = 8'h29;
  picture_data[ 3447 ] = 8'h23;
  picture_data[ 3448 ] = 8'h39;
  picture_data[ 3449 ] = 8'hC5;
  picture_data[ 3450 ] = 8'h39;
  picture_data[ 3451 ] = 8'hE5;
  picture_data[ 3452 ] = 8'h31;
  picture_data[ 3453 ] = 8'h83;
  picture_data[ 3454 ] = 8'h21;
  picture_data[ 3455 ] = 8'h22;
  picture_data[ 3456 ] = 8'h21;
  picture_data[ 3457 ] = 8'h22;
  picture_data[ 3458 ] = 8'h31;
  picture_data[ 3459 ] = 8'hA4;
  picture_data[ 3460 ] = 8'h41;
  picture_data[ 3461 ] = 8'hE5;
  picture_data[ 3462 ] = 8'h41;
  picture_data[ 3463 ] = 8'hC5;
  picture_data[ 3464 ] = 8'h39;
  picture_data[ 3465 ] = 8'hC4;
  picture_data[ 3466 ] = 8'h39;
  picture_data[ 3467 ] = 8'hA3;
  picture_data[ 3468 ] = 8'h41;
  picture_data[ 3469 ] = 8'hC3;
  picture_data[ 3470 ] = 8'h52;
  picture_data[ 3471 ] = 8'h24;
  picture_data[ 3472 ] = 8'h72;
  picture_data[ 3473 ] = 8'hC6;
  picture_data[ 3474 ] = 8'h7A;
  picture_data[ 3475 ] = 8'hE6;
  picture_data[ 3476 ] = 8'h7A;
  picture_data[ 3477 ] = 8'h85;
  picture_data[ 3478 ] = 8'h8B;
  picture_data[ 3479 ] = 8'h27;
  picture_data[ 3480 ] = 8'h6A;
  picture_data[ 3481 ] = 8'h24;
  picture_data[ 3482 ] = 8'h62;
  picture_data[ 3483 ] = 8'h23;
  picture_data[ 3484 ] = 8'hB4;
  picture_data[ 3485 ] = 8'hCE;
  picture_data[ 3486 ] = 8'hB5;
  picture_data[ 3487 ] = 8'h2F;
  picture_data[ 3488 ] = 8'hAD;
  picture_data[ 3489 ] = 8'h2F;
  picture_data[ 3490 ] = 8'hAC;
  picture_data[ 3491 ] = 8'hEF;
  picture_data[ 3492 ] = 8'hC5;
  picture_data[ 3493 ] = 8'h92;
  picture_data[ 3494 ] = 8'hEE;
  picture_data[ 3495 ] = 8'hB7;
  picture_data[ 3496 ] = 8'h08;
  picture_data[ 3497 ] = 8'hA2;
  picture_data[ 3498 ] = 8'h00;
  picture_data[ 3499 ] = 8'hA2;
  picture_data[ 3500 ] = 8'h08;
  picture_data[ 3501 ] = 8'hE3;
  picture_data[ 3502 ] = 8'h11;
  picture_data[ 3503 ] = 8'h24;
  picture_data[ 3504 ] = 8'h11;
  picture_data[ 3505 ] = 8'h24;
  picture_data[ 3506 ] = 8'h10;
  picture_data[ 3507 ] = 8'hE4;
  picture_data[ 3508 ] = 8'h10;
  picture_data[ 3509 ] = 8'hC3;
  picture_data[ 3510 ] = 8'h10;
  picture_data[ 3511 ] = 8'hE3;
  picture_data[ 3512 ] = 8'h21;
  picture_data[ 3513 ] = 8'h64;
  picture_data[ 3514 ] = 8'h29;
  picture_data[ 3515 ] = 8'hA5;
  picture_data[ 3516 ] = 8'h19;
  picture_data[ 3517 ] = 8'h63;
  picture_data[ 3518 ] = 8'h21;
  picture_data[ 3519 ] = 8'h83;
  picture_data[ 3520 ] = 8'h29;
  picture_data[ 3521 ] = 8'hE5;
  picture_data[ 3522 ] = 8'h21;
  picture_data[ 3523 ] = 8'h63;
  picture_data[ 3524 ] = 8'h29;
  picture_data[ 3525 ] = 8'h84;
  picture_data[ 3526 ] = 8'h5A;
  picture_data[ 3527 ] = 8'hA8;
  picture_data[ 3528 ] = 8'h5A;
  picture_data[ 3529 ] = 8'hC8;
  picture_data[ 3530 ] = 8'h52;
  picture_data[ 3531 ] = 8'h67;
  picture_data[ 3532 ] = 8'h6A;
  picture_data[ 3533 ] = 8'hEA;
  picture_data[ 3534 ] = 8'h7B;
  picture_data[ 3535 ] = 8'h2B;
  picture_data[ 3536 ] = 8'h72;
  picture_data[ 3537 ] = 8'hA8;
  picture_data[ 3538 ] = 8'h72;
  picture_data[ 3539 ] = 8'hA7;
  picture_data[ 3540 ] = 8'h62;
  picture_data[ 3541 ] = 8'h67;
  picture_data[ 3542 ] = 8'h6A;
  picture_data[ 3543 ] = 8'hA9;
  picture_data[ 3544 ] = 8'h6A;
  picture_data[ 3545 ] = 8'hAA;
  picture_data[ 3546 ] = 8'h51;
  picture_data[ 3547 ] = 8'hC7;
  picture_data[ 3548 ] = 8'h6A;
  picture_data[ 3549 ] = 8'hAA;
  picture_data[ 3550 ] = 8'h7B;
  picture_data[ 3551 ] = 8'h2B;
  picture_data[ 3552 ] = 8'h73;
  picture_data[ 3553 ] = 8'h2B;
  picture_data[ 3554 ] = 8'h28;
  picture_data[ 3555 ] = 8'hC3;
  picture_data[ 3556 ] = 8'h29;
  picture_data[ 3557 ] = 8'h03;
  picture_data[ 3558 ] = 8'h31;
  picture_data[ 3559 ] = 8'h65;
  picture_data[ 3560 ] = 8'h28;
  picture_data[ 3561 ] = 8'hE3;
  picture_data[ 3562 ] = 8'h31;
  picture_data[ 3563 ] = 8'h45;
  picture_data[ 3564 ] = 8'h31;
  picture_data[ 3565 ] = 8'h65;
  picture_data[ 3566 ] = 8'h29;
  picture_data[ 3567 ] = 8'h24;
  picture_data[ 3568 ] = 8'h39;
  picture_data[ 3569 ] = 8'h86;
  picture_data[ 3570 ] = 8'h31;
  picture_data[ 3571 ] = 8'h65;
  picture_data[ 3572 ] = 8'h29;
  picture_data[ 3573 ] = 8'h05;
  picture_data[ 3574 ] = 8'h31;
  picture_data[ 3575 ] = 8'h25;
  picture_data[ 3576 ] = 8'h39;
  picture_data[ 3577 ] = 8'h87;
  picture_data[ 3578 ] = 8'h5A;
  picture_data[ 3579 ] = 8'h8A;
  picture_data[ 3580 ] = 8'h39;
  picture_data[ 3581 ] = 8'h65;
  picture_data[ 3582 ] = 8'h52;
  picture_data[ 3583 ] = 8'h07;
  picture_data[ 3584 ] = 8'h49;
  picture_data[ 3585 ] = 8'hC6;
  picture_data[ 3586 ] = 8'h51;
  picture_data[ 3587 ] = 8'hE6;
  picture_data[ 3588 ] = 8'h49;
  picture_data[ 3589 ] = 8'hC6;
  picture_data[ 3590 ] = 8'h39;
  picture_data[ 3591 ] = 8'h64;
  picture_data[ 3592 ] = 8'h5A;
  picture_data[ 3593 ] = 8'h89;
  picture_data[ 3594 ] = 8'h31;
  picture_data[ 3595 ] = 8'h85;
  picture_data[ 3596 ] = 8'h4A;
  picture_data[ 3597 ] = 8'h27;
  picture_data[ 3598 ] = 8'h21;
  picture_data[ 3599 ] = 8'h02;
  picture_data[ 3600 ] = 8'h31;
  picture_data[ 3601 ] = 8'h63;
  picture_data[ 3602 ] = 8'h39;
  picture_data[ 3603 ] = 8'hA4;
  picture_data[ 3604 ] = 8'h31;
  picture_data[ 3605 ] = 8'hC4;
  picture_data[ 3606 ] = 8'h29;
  picture_data[ 3607 ] = 8'h83;
  picture_data[ 3608 ] = 8'h42;
  picture_data[ 3609 ] = 8'h06;
  picture_data[ 3610 ] = 8'h42;
  picture_data[ 3611 ] = 8'h06;
  picture_data[ 3612 ] = 8'h39;
  picture_data[ 3613 ] = 8'hA4;
  picture_data[ 3614 ] = 8'h31;
  picture_data[ 3615 ] = 8'hA4;
  picture_data[ 3616 ] = 8'h39;
  picture_data[ 3617 ] = 8'hC4;
  picture_data[ 3618 ] = 8'h41;
  picture_data[ 3619 ] = 8'hE4;
  picture_data[ 3620 ] = 8'h39;
  picture_data[ 3621 ] = 8'hA3;
  picture_data[ 3622 ] = 8'h41;
  picture_data[ 3623 ] = 8'hC3;
  picture_data[ 3624 ] = 8'h49;
  picture_data[ 3625 ] = 8'hC3;
  picture_data[ 3626 ] = 8'h62;
  picture_data[ 3627 ] = 8'h44;
  picture_data[ 3628 ] = 8'h6A;
  picture_data[ 3629 ] = 8'h44;
  picture_data[ 3630 ] = 8'h59;
  picture_data[ 3631 ] = 8'hE3;
  picture_data[ 3632 ] = 8'h62;
  picture_data[ 3633 ] = 8'h03;
  picture_data[ 3634 ] = 8'h6A;
  picture_data[ 3635 ] = 8'h44;
  picture_data[ 3636 ] = 8'hB4;
  picture_data[ 3637 ] = 8'hCE;
  picture_data[ 3638 ] = 8'hB5;
  picture_data[ 3639 ] = 8'h0F;
  picture_data[ 3640 ] = 8'hAD;
  picture_data[ 3641 ] = 8'h0F;
  picture_data[ 3642 ] = 8'hAC;
  picture_data[ 3643 ] = 8'hEF;
  picture_data[ 3644 ] = 8'hC5;
  picture_data[ 3645 ] = 8'h72;
  picture_data[ 3646 ] = 8'hEE;
  picture_data[ 3647 ] = 8'h97;
  picture_data[ 3648 ] = 8'h21;
  picture_data[ 3649 ] = 8'h86;
  picture_data[ 3650 ] = 8'h19;
  picture_data[ 3651 ] = 8'h65;
  picture_data[ 3652 ] = 8'h08;
  picture_data[ 3653 ] = 8'hE3;
  picture_data[ 3654 ] = 8'h11;
  picture_data[ 3655 ] = 8'h24;
  picture_data[ 3656 ] = 8'h08;
  picture_data[ 3657 ] = 8'hE4;
  picture_data[ 3658 ] = 8'h08;
  picture_data[ 3659 ] = 8'hE4;
  picture_data[ 3660 ] = 8'h10;
  picture_data[ 3661 ] = 8'hE4;
  picture_data[ 3662 ] = 8'h10;
  picture_data[ 3663 ] = 8'hC3;
  picture_data[ 3664 ] = 8'h29;
  picture_data[ 3665 ] = 8'hA6;
  picture_data[ 3666 ] = 8'h29;
  picture_data[ 3667 ] = 8'hA5;
  picture_data[ 3668 ] = 8'h19;
  picture_data[ 3669 ] = 8'h42;
  picture_data[ 3670 ] = 8'h29;
  picture_data[ 3671 ] = 8'hA3;
  picture_data[ 3672 ] = 8'h19;
  picture_data[ 3673 ] = 8'h42;
  picture_data[ 3674 ] = 8'h19;
  picture_data[ 3675 ] = 8'h01;
  picture_data[ 3676 ] = 8'h29;
  picture_data[ 3677 ] = 8'h84;
  picture_data[ 3678 ] = 8'h52;
  picture_data[ 3679 ] = 8'hA8;
  picture_data[ 3680 ] = 8'h52;
  picture_data[ 3681 ] = 8'h86;
  picture_data[ 3682 ] = 8'h52;
  picture_data[ 3683 ] = 8'h66;
  picture_data[ 3684 ] = 8'h5A;
  picture_data[ 3685 ] = 8'h67;
  picture_data[ 3686 ] = 8'h51;
  picture_data[ 3687 ] = 8'hC5;
  picture_data[ 3688 ] = 8'h5A;
  picture_data[ 3689 ] = 8'h05;
  picture_data[ 3690 ] = 8'h72;
  picture_data[ 3691 ] = 8'hA8;
  picture_data[ 3692 ] = 8'h6A;
  picture_data[ 3693 ] = 8'hA8;
  picture_data[ 3694 ] = 8'h62;
  picture_data[ 3695 ] = 8'h68;
  picture_data[ 3696 ] = 8'h5A;
  picture_data[ 3697 ] = 8'h48;
  picture_data[ 3698 ] = 8'h5A;
  picture_data[ 3699 ] = 8'h68;
  picture_data[ 3700 ] = 8'h62;
  picture_data[ 3701 ] = 8'h69;
  picture_data[ 3702 ] = 8'h41;
  picture_data[ 3703 ] = 8'h64;
  picture_data[ 3704 ] = 8'h39;
  picture_data[ 3705 ] = 8'h44;
  picture_data[ 3706 ] = 8'h28;
  picture_data[ 3707 ] = 8'hE2;
  picture_data[ 3708 ] = 8'h31;
  picture_data[ 3709 ] = 8'h44;
  picture_data[ 3710 ] = 8'h29;
  picture_data[ 3711 ] = 8'h04;
  picture_data[ 3712 ] = 8'h28;
  picture_data[ 3713 ] = 8'hE3;
  picture_data[ 3714 ] = 8'h28;
  picture_data[ 3715 ] = 8'hE3;
  picture_data[ 3716 ] = 8'h20;
  picture_data[ 3717 ] = 8'hA2;
  picture_data[ 3718 ] = 8'h39;
  picture_data[ 3719 ] = 8'h85;
  picture_data[ 3720 ] = 8'h39;
  picture_data[ 3721 ] = 8'hA6;
  picture_data[ 3722 ] = 8'h41;
  picture_data[ 3723 ] = 8'hE8;
  picture_data[ 3724 ] = 8'h39;
  picture_data[ 3725 ] = 8'h87;
  picture_data[ 3726 ] = 8'h39;
  picture_data[ 3727 ] = 8'h87;
  picture_data[ 3728 ] = 8'h20;
  picture_data[ 3729 ] = 8'hC4;
  picture_data[ 3730 ] = 8'h5A;
  picture_data[ 3731 ] = 8'h8B;
  picture_data[ 3732 ] = 8'h41;
  picture_data[ 3733 ] = 8'hC7;
  picture_data[ 3734 ] = 8'h49;
  picture_data[ 3735 ] = 8'hE7;
  picture_data[ 3736 ] = 8'h52;
  picture_data[ 3737 ] = 8'h07;
  picture_data[ 3738 ] = 8'h49;
  picture_data[ 3739 ] = 8'hC6;
  picture_data[ 3740 ] = 8'h39;
  picture_data[ 3741 ] = 8'h44;
  picture_data[ 3742 ] = 8'h41;
  picture_data[ 3743 ] = 8'hC6;
  picture_data[ 3744 ] = 8'h39;
  picture_data[ 3745 ] = 8'h85;
  picture_data[ 3746 ] = 8'h21;
  picture_data[ 3747 ] = 8'h23;
  picture_data[ 3748 ] = 8'h29;
  picture_data[ 3749 ] = 8'h43;
  picture_data[ 3750 ] = 8'h29;
  picture_data[ 3751 ] = 8'h43;
  picture_data[ 3752 ] = 8'h21;
  picture_data[ 3753 ] = 8'h02;
  picture_data[ 3754 ] = 8'h39;
  picture_data[ 3755 ] = 8'hE5;
  picture_data[ 3756 ] = 8'h29;
  picture_data[ 3757 ] = 8'h63;
  picture_data[ 3758 ] = 8'h21;
  picture_data[ 3759 ] = 8'h42;
  picture_data[ 3760 ] = 8'h31;
  picture_data[ 3761 ] = 8'hC4;
  picture_data[ 3762 ] = 8'h31;
  picture_data[ 3763 ] = 8'hC4;
  picture_data[ 3764 ] = 8'h42;
  picture_data[ 3765 ] = 8'h25;
  picture_data[ 3766 ] = 8'h39;
  picture_data[ 3767 ] = 8'hE4;
  picture_data[ 3768 ] = 8'h42;
  picture_data[ 3769 ] = 8'h05;
  picture_data[ 3770 ] = 8'h42;
  picture_data[ 3771 ] = 8'h04;
  picture_data[ 3772 ] = 8'h4A;
  picture_data[ 3773 ] = 8'h45;
  picture_data[ 3774 ] = 8'h6B;
  picture_data[ 3775 ] = 8'h29;
  picture_data[ 3776 ] = 8'h5A;
  picture_data[ 3777 ] = 8'h46;
  picture_data[ 3778 ] = 8'h62;
  picture_data[ 3779 ] = 8'h66;
  picture_data[ 3780 ] = 8'h5A;
  picture_data[ 3781 ] = 8'h05;
  picture_data[ 3782 ] = 8'h59;
  picture_data[ 3783 ] = 8'hE4;
  picture_data[ 3784 ] = 8'h62;
  picture_data[ 3785 ] = 8'h04;
  picture_data[ 3786 ] = 8'h72;
  picture_data[ 3787 ] = 8'h66;
  picture_data[ 3788 ] = 8'hBC;
  picture_data[ 3789 ] = 8'hEF;
  picture_data[ 3790 ] = 8'hB4;
  picture_data[ 3791 ] = 8'hCF;
  picture_data[ 3792 ] = 8'hB4;
  picture_data[ 3793 ] = 8'hEF;
  picture_data[ 3794 ] = 8'hAC;
  picture_data[ 3795 ] = 8'hCF;
  picture_data[ 3796 ] = 8'hBD;
  picture_data[ 3797 ] = 8'h51;
  picture_data[ 3798 ] = 8'hEE;
  picture_data[ 3799 ] = 8'hB7;
  picture_data[ 3800 ] = 8'h4A;
  picture_data[ 3801 ] = 8'hCA;
  picture_data[ 3802 ] = 8'h08;
  picture_data[ 3803 ] = 8'hC2;
  picture_data[ 3804 ] = 8'h11;
  picture_data[ 3805 ] = 8'h24;
  picture_data[ 3806 ] = 8'h11;
  picture_data[ 3807 ] = 8'h24;
  picture_data[ 3808 ] = 8'h08;
  picture_data[ 3809 ] = 8'hE3;
  picture_data[ 3810 ] = 8'h00;
  picture_data[ 3811 ] = 8'hA2;
  picture_data[ 3812 ] = 8'h10;
  picture_data[ 3813 ] = 8'hC3;
  picture_data[ 3814 ] = 8'h29;
  picture_data[ 3815 ] = 8'h86;
  picture_data[ 3816 ] = 8'h29;
  picture_data[ 3817 ] = 8'h86;
  picture_data[ 3818 ] = 8'h19;
  picture_data[ 3819 ] = 8'h03;
  picture_data[ 3820 ] = 8'h21;
  picture_data[ 3821 ] = 8'h84;
  picture_data[ 3822 ] = 8'h29;
  picture_data[ 3823 ] = 8'hC4;
  picture_data[ 3824 ] = 8'h29;
  picture_data[ 3825 ] = 8'hA3;
  picture_data[ 3826 ] = 8'h19;
  picture_data[ 3827 ] = 8'h01;
  picture_data[ 3828 ] = 8'h4A;
  picture_data[ 3829 ] = 8'h47;
  picture_data[ 3830 ] = 8'h5A;
  picture_data[ 3831 ] = 8'hC9;
  picture_data[ 3832 ] = 8'h42;
  picture_data[ 3833 ] = 8'h45;
  picture_data[ 3834 ] = 8'h39;
  picture_data[ 3835 ] = 8'hC3;
  picture_data[ 3836 ] = 8'h39;
  picture_data[ 3837 ] = 8'h63;
  picture_data[ 3838 ] = 8'h5A;
  picture_data[ 3839 ] = 8'h47;
  picture_data[ 3840 ] = 8'h51;
  picture_data[ 3841 ] = 8'hE5;
  picture_data[ 3842 ] = 8'h5A;
  picture_data[ 3843 ] = 8'h26;
  picture_data[ 3844 ] = 8'h5A;
  picture_data[ 3845 ] = 8'h87;
  picture_data[ 3846 ] = 8'h62;
  picture_data[ 3847 ] = 8'h88;
  picture_data[ 3848 ] = 8'h41;
  picture_data[ 3849 ] = 8'hE5;
  picture_data[ 3850 ] = 8'h41;
  picture_data[ 3851 ] = 8'hC5;
  picture_data[ 3852 ] = 8'h39;
  picture_data[ 3853 ] = 8'h84;
  picture_data[ 3854 ] = 8'h31;
  picture_data[ 3855 ] = 8'h23;
  picture_data[ 3856 ] = 8'h31;
  picture_data[ 3857 ] = 8'h24;
  picture_data[ 3858 ] = 8'h20;
  picture_data[ 3859 ] = 8'hC2;
  picture_data[ 3860 ] = 8'h29;
  picture_data[ 3861 ] = 8'h03;
  picture_data[ 3862 ] = 8'h28;
  picture_data[ 3863 ] = 8'hE3;
  picture_data[ 3864 ] = 8'h20;
  picture_data[ 3865 ] = 8'h82;
  picture_data[ 3866 ] = 8'h20;
  picture_data[ 3867 ] = 8'hA2;
  picture_data[ 3868 ] = 8'h20;
  picture_data[ 3869 ] = 8'hC2;
  picture_data[ 3870 ] = 8'h39;
  picture_data[ 3871 ] = 8'h65;
  picture_data[ 3872 ] = 8'h5A;
  picture_data[ 3873 ] = 8'h69;
  picture_data[ 3874 ] = 8'h39;
  picture_data[ 3875 ] = 8'h86;
  picture_data[ 3876 ] = 8'h21;
  picture_data[ 3877 ] = 8'h04;
  picture_data[ 3878 ] = 8'h31;
  picture_data[ 3879 ] = 8'h66;
  picture_data[ 3880 ] = 8'h18;
  picture_data[ 3881 ] = 8'hA3;
  picture_data[ 3882 ] = 8'h41;
  picture_data[ 3883 ] = 8'hE8;
  picture_data[ 3884 ] = 8'h39;
  picture_data[ 3885 ] = 8'h86;
  picture_data[ 3886 ] = 8'h41;
  picture_data[ 3887 ] = 8'hA6;
  picture_data[ 3888 ] = 8'h5A;
  picture_data[ 3889 ] = 8'h68;
  picture_data[ 3890 ] = 8'h41;
  picture_data[ 3891 ] = 8'h85;
  picture_data[ 3892 ] = 8'h28;
  picture_data[ 3893 ] = 8'hC2;
  picture_data[ 3894 ] = 8'h41;
  picture_data[ 3895 ] = 8'hA5;
  picture_data[ 3896 ] = 8'h29;
  picture_data[ 3897 ] = 8'h44;
  picture_data[ 3898 ] = 8'h21;
  picture_data[ 3899 ] = 8'h23;
  picture_data[ 3900 ] = 8'h31;
  picture_data[ 3901 ] = 8'h84;
  picture_data[ 3902 ] = 8'h31;
  picture_data[ 3903 ] = 8'hA4;
  picture_data[ 3904 ] = 8'h21;
  picture_data[ 3905 ] = 8'h02;
  picture_data[ 3906 ] = 8'h29;
  picture_data[ 3907 ] = 8'h63;
  picture_data[ 3908 ] = 8'h21;
  picture_data[ 3909 ] = 8'h43;
  picture_data[ 3910 ] = 8'h29;
  picture_data[ 3911 ] = 8'h83;
  picture_data[ 3912 ] = 8'h39;
  picture_data[ 3913 ] = 8'hC4;
  picture_data[ 3914 ] = 8'h31;
  picture_data[ 3915 ] = 8'hC4;
  picture_data[ 3916 ] = 8'h39;
  picture_data[ 3917 ] = 8'hE4;
  picture_data[ 3918 ] = 8'h39;
  picture_data[ 3919 ] = 8'hE4;
  picture_data[ 3920 ] = 8'h39;
  picture_data[ 3921 ] = 8'hC4;
  picture_data[ 3922 ] = 8'h39;
  picture_data[ 3923 ] = 8'hC3;
  picture_data[ 3924 ] = 8'h42;
  picture_data[ 3925 ] = 8'h04;
  picture_data[ 3926 ] = 8'h41;
  picture_data[ 3927 ] = 8'hE4;
  picture_data[ 3928 ] = 8'h7B;
  picture_data[ 3929 ] = 8'h4A;
  picture_data[ 3930 ] = 8'h6A;
  picture_data[ 3931 ] = 8'hA8;
  picture_data[ 3932 ] = 8'h62;
  picture_data[ 3933 ] = 8'h46;
  picture_data[ 3934 ] = 8'h49;
  picture_data[ 3935 ] = 8'hA3;
  picture_data[ 3936 ] = 8'h51;
  picture_data[ 3937 ] = 8'hA3;
  picture_data[ 3938 ] = 8'h62;
  picture_data[ 3939 ] = 8'h25;
  picture_data[ 3940 ] = 8'hA4;
  picture_data[ 3941 ] = 8'h0C;
  picture_data[ 3942 ] = 8'hB4;
  picture_data[ 3943 ] = 8'hCF;
  picture_data[ 3944 ] = 8'hAC;
  picture_data[ 3945 ] = 8'hAE;
  picture_data[ 3946 ] = 8'hAC;
  picture_data[ 3947 ] = 8'hCF;
  picture_data[ 3948 ] = 8'hB4;
  picture_data[ 3949 ] = 8'hF0;
  picture_data[ 3950 ] = 8'hDE;
  picture_data[ 3951 ] = 8'h55;
  picture_data[ 3952 ] = 8'h5B;
  picture_data[ 3953 ] = 8'h4B;
  picture_data[ 3954 ] = 8'h10;
  picture_data[ 3955 ] = 8'hE1;
  picture_data[ 3956 ] = 8'h00;
  picture_data[ 3957 ] = 8'hA1;
  picture_data[ 3958 ] = 8'h08;
  picture_data[ 3959 ] = 8'hC3;
  picture_data[ 3960 ] = 8'h08;
  picture_data[ 3961 ] = 8'hA2;
  picture_data[ 3962 ] = 8'h19;
  picture_data[ 3963 ] = 8'h24;
  picture_data[ 3964 ] = 8'h21;
  picture_data[ 3965 ] = 8'h45;
  picture_data[ 3966 ] = 8'h29;
  picture_data[ 3967 ] = 8'h66;
  picture_data[ 3968 ] = 8'h10;
  picture_data[ 3969 ] = 8'hA2;
  picture_data[ 3970 ] = 8'h31;
  picture_data[ 3971 ] = 8'hA6;
  picture_data[ 3972 ] = 8'h31;
  picture_data[ 3973 ] = 8'hE6;
  picture_data[ 3974 ] = 8'h31;
  picture_data[ 3975 ] = 8'hC5;
  picture_data[ 3976 ] = 8'h19;
  picture_data[ 3977 ] = 8'h22;
  picture_data[ 3978 ] = 8'h29;
  picture_data[ 3979 ] = 8'h83;
  picture_data[ 3980 ] = 8'h42;
  picture_data[ 3981 ] = 8'h06;
  picture_data[ 3982 ] = 8'h4A;
  picture_data[ 3983 ] = 8'h67;
  picture_data[ 3984 ] = 8'h39;
  picture_data[ 3985 ] = 8'hE5;
  picture_data[ 3986 ] = 8'h39;
  picture_data[ 3987 ] = 8'hC4;
  picture_data[ 3988 ] = 8'h31;
  picture_data[ 3989 ] = 8'h83;
  picture_data[ 3990 ] = 8'h52;
  picture_data[ 3991 ] = 8'h47;
  picture_data[ 3992 ] = 8'h41;
  picture_data[ 3993 ] = 8'hA4;
  picture_data[ 3994 ] = 8'h52;
  picture_data[ 3995 ] = 8'h26;
  picture_data[ 3996 ] = 8'h52;
  picture_data[ 3997 ] = 8'h67;
  picture_data[ 3998 ] = 8'h39;
  picture_data[ 3999 ] = 8'h83;
  picture_data[ 4000 ] = 8'h29;
  picture_data[ 4001 ] = 8'h42;
  picture_data[ 4002 ] = 8'h29;
  picture_data[ 4003 ] = 8'h21;
  picture_data[ 4004 ] = 8'h31;
  picture_data[ 4005 ] = 8'h63;
  picture_data[ 4006 ] = 8'h39;
  picture_data[ 4007 ] = 8'h64;
  picture_data[ 4008 ] = 8'h20;
  picture_data[ 4009 ] = 8'hC2;
  picture_data[ 4010 ] = 8'h20;
  picture_data[ 4011 ] = 8'hE3;
  picture_data[ 4012 ] = 8'h29;
  picture_data[ 4013 ] = 8'h03;
  picture_data[ 4014 ] = 8'h18;
  picture_data[ 4015 ] = 8'hA1;
  picture_data[ 4016 ] = 8'h28;
  picture_data[ 4017 ] = 8'hE3;
  picture_data[ 4018 ] = 8'h39;
  picture_data[ 4019 ] = 8'h86;
  picture_data[ 4020 ] = 8'h39;
  picture_data[ 4021 ] = 8'h65;
  picture_data[ 4022 ] = 8'h29;
  picture_data[ 4023 ] = 8'h23;
  picture_data[ 4024 ] = 8'h39;
  picture_data[ 4025 ] = 8'h65;
  picture_data[ 4026 ] = 8'h4A;
  picture_data[ 4027 ] = 8'h08;
  picture_data[ 4028 ] = 8'h4A;
  picture_data[ 4029 ] = 8'h49;
  picture_data[ 4030 ] = 8'h52;
  picture_data[ 4031 ] = 8'h4A;
  picture_data[ 4032 ] = 8'h29;
  picture_data[ 4033 ] = 8'h05;
  picture_data[ 4034 ] = 8'h29;
  picture_data[ 4035 ] = 8'h25;
  picture_data[ 4036 ] = 8'h39;
  picture_data[ 4037 ] = 8'h85;
  picture_data[ 4038 ] = 8'h4A;
  picture_data[ 4039 ] = 8'h07;
  picture_data[ 4040 ] = 8'h49;
  picture_data[ 4041 ] = 8'hE6;
  picture_data[ 4042 ] = 8'h41;
  picture_data[ 4043 ] = 8'hA5;
  picture_data[ 4044 ] = 8'h39;
  picture_data[ 4045 ] = 8'h65;
  picture_data[ 4046 ] = 8'h39;
  picture_data[ 4047 ] = 8'h65;
  picture_data[ 4048 ] = 8'h4A;
  picture_data[ 4049 ] = 8'h28;
  picture_data[ 4050 ] = 8'h29;
  picture_data[ 4051 ] = 8'h85;
  picture_data[ 4052 ] = 8'h21;
  picture_data[ 4053 ] = 8'h02;
  picture_data[ 4054 ] = 8'h21;
  picture_data[ 4055 ] = 8'h23;
  picture_data[ 4056 ] = 8'h18;
  picture_data[ 4057 ] = 8'hE1;
  picture_data[ 4058 ] = 8'h21;
  picture_data[ 4059 ] = 8'h02;
  picture_data[ 4060 ] = 8'h29;
  picture_data[ 4061 ] = 8'h63;
  picture_data[ 4062 ] = 8'h4A;
  picture_data[ 4063 ] = 8'h46;
  picture_data[ 4064 ] = 8'h4A;
  picture_data[ 4065 ] = 8'h66;
  picture_data[ 4066 ] = 8'h42;
  picture_data[ 4067 ] = 8'h25;
  picture_data[ 4068 ] = 8'h39;
  picture_data[ 4069 ] = 8'hE4;
  picture_data[ 4070 ] = 8'h31;
  picture_data[ 4071 ] = 8'hC3;
  picture_data[ 4072 ] = 8'h31;
  picture_data[ 4073 ] = 8'hA3;
  picture_data[ 4074 ] = 8'h39;
  picture_data[ 4075 ] = 8'hE4;
  picture_data[ 4076 ] = 8'h39;
  picture_data[ 4077 ] = 8'hE4;
  picture_data[ 4078 ] = 8'h42;
  picture_data[ 4079 ] = 8'h04;
  picture_data[ 4080 ] = 8'h62;
  picture_data[ 4081 ] = 8'hC8;
  picture_data[ 4082 ] = 8'h52;
  picture_data[ 4083 ] = 8'h66;
  picture_data[ 4084 ] = 8'h49;
  picture_data[ 4085 ] = 8'hE4;
  picture_data[ 4086 ] = 8'h39;
  picture_data[ 4087 ] = 8'h62;
  picture_data[ 4088 ] = 8'h41;
  picture_data[ 4089 ] = 8'h82;
  picture_data[ 4090 ] = 8'h51;
  picture_data[ 4091 ] = 8'hE3;
  picture_data[ 4092 ] = 8'hA4;
  picture_data[ 4093 ] = 8'h4D;
  picture_data[ 4094 ] = 8'hB4;
  picture_data[ 4095 ] = 8'hEF;
  picture_data[ 4096 ] = 8'hB4;
  picture_data[ 4097 ] = 8'hCF;
  picture_data[ 4098 ] = 8'hAC;
  picture_data[ 4099 ] = 8'hD0;
  picture_data[ 4100 ] = 8'hBD;
  picture_data[ 4101 ] = 8'h72;
  picture_data[ 4102 ] = 8'hC5;
  picture_data[ 4103 ] = 8'hD4;
  picture_data[ 4104 ] = 8'h4A;
  picture_data[ 4105 ] = 8'hA8;
  picture_data[ 4106 ] = 8'h42;
  picture_data[ 4107 ] = 8'h67;
  picture_data[ 4108 ] = 8'h00;
  picture_data[ 4109 ] = 8'h20;
  picture_data[ 4110 ] = 8'h08;
  picture_data[ 4111 ] = 8'hE2;
  picture_data[ 4112 ] = 8'h11;
  picture_data[ 4113 ] = 8'h03;
  picture_data[ 4114 ] = 8'h29;
  picture_data[ 4115 ] = 8'hA6;
  picture_data[ 4116 ] = 8'h21;
  picture_data[ 4117 ] = 8'h65;
  picture_data[ 4118 ] = 8'h10;
  picture_data[ 4119 ] = 8'hE3;
  picture_data[ 4120 ] = 8'h18;
  picture_data[ 4121 ] = 8'hE3;
  picture_data[ 4122 ] = 8'h21;
  picture_data[ 4123 ] = 8'h24;
  picture_data[ 4124 ] = 8'h29;
  picture_data[ 4125 ] = 8'h85;
  picture_data[ 4126 ] = 8'h21;
  picture_data[ 4127 ] = 8'h84;
  picture_data[ 4128 ] = 8'h10;
  picture_data[ 4129 ] = 8'hE1;
  picture_data[ 4130 ] = 8'h10;
  picture_data[ 4131 ] = 8'hC1;
  picture_data[ 4132 ] = 8'h31;
  picture_data[ 4133 ] = 8'h85;
  picture_data[ 4134 ] = 8'h31;
  picture_data[ 4135 ] = 8'h85;
  picture_data[ 4136 ] = 8'h31;
  picture_data[ 4137 ] = 8'h84;
  picture_data[ 4138 ] = 8'h18;
  picture_data[ 4139 ] = 8'hC0;
  picture_data[ 4140 ] = 8'h42;
  picture_data[ 4141 ] = 8'h05;
  picture_data[ 4142 ] = 8'h31;
  picture_data[ 4143 ] = 8'h63;
  picture_data[ 4144 ] = 8'h21;
  picture_data[ 4145 ] = 8'h22;
  picture_data[ 4146 ] = 8'h4A;
  picture_data[ 4147 ] = 8'h26;
  picture_data[ 4148 ] = 8'h10;
  picture_data[ 4149 ] = 8'h80;
  picture_data[ 4150 ] = 8'h18;
  picture_data[ 4151 ] = 8'hC0;
  picture_data[ 4152 ] = 8'h29;
  picture_data[ 4153 ] = 8'h62;
  picture_data[ 4154 ] = 8'h31;
  picture_data[ 4155 ] = 8'h62;
  picture_data[ 4156 ] = 8'h31;
  picture_data[ 4157 ] = 8'h63;
  picture_data[ 4158 ] = 8'h31;
  picture_data[ 4159 ] = 8'h43;
  picture_data[ 4160 ] = 8'h29;
  picture_data[ 4161 ] = 8'h03;
  picture_data[ 4162 ] = 8'h20;
  picture_data[ 4163 ] = 8'hC2;
  picture_data[ 4164 ] = 8'h10;
  picture_data[ 4165 ] = 8'h60;
  picture_data[ 4166 ] = 8'h39;
  picture_data[ 4167 ] = 8'h65;
  picture_data[ 4168 ] = 8'h31;
  picture_data[ 4169 ] = 8'h44;
  picture_data[ 4170 ] = 8'h20;
  picture_data[ 4171 ] = 8'hA2;
  picture_data[ 4172 ] = 8'h31;
  picture_data[ 4173 ] = 8'h44;
  picture_data[ 4174 ] = 8'h31;
  picture_data[ 4175 ] = 8'h44;
  picture_data[ 4176 ] = 8'h31;
  picture_data[ 4177 ] = 8'h44;
  picture_data[ 4178 ] = 8'h29;
  picture_data[ 4179 ] = 8'h24;
  picture_data[ 4180 ] = 8'h41;
  picture_data[ 4181 ] = 8'hE7;
  picture_data[ 4182 ] = 8'h41;
  picture_data[ 4183 ] = 8'hE7;
  picture_data[ 4184 ] = 8'h31;
  picture_data[ 4185 ] = 8'h45;
  picture_data[ 4186 ] = 8'h18;
  picture_data[ 4187 ] = 8'hA2;
  picture_data[ 4188 ] = 8'h39;
  picture_data[ 4189 ] = 8'h85;
  picture_data[ 4190 ] = 8'h41;
  picture_data[ 4191 ] = 8'hE6;
  picture_data[ 4192 ] = 8'h39;
  picture_data[ 4193 ] = 8'h84;
  picture_data[ 4194 ] = 8'h4A;
  picture_data[ 4195 ] = 8'h06;
  picture_data[ 4196 ] = 8'h62;
  picture_data[ 4197 ] = 8'hA9;
  picture_data[ 4198 ] = 8'h39;
  picture_data[ 4199 ] = 8'hA5;
  picture_data[ 4200 ] = 8'h42;
  picture_data[ 4201 ] = 8'h07;
  picture_data[ 4202 ] = 8'h31;
  picture_data[ 4203 ] = 8'hA5;
  picture_data[ 4204 ] = 8'h21;
  picture_data[ 4205 ] = 8'h43;
  picture_data[ 4206 ] = 8'h29;
  picture_data[ 4207 ] = 8'h84;
  picture_data[ 4208 ] = 8'h29;
  picture_data[ 4209 ] = 8'h64;
  picture_data[ 4210 ] = 8'h21;
  picture_data[ 4211 ] = 8'h23;
  picture_data[ 4212 ] = 8'h21;
  picture_data[ 4213 ] = 8'h02;
  picture_data[ 4214 ] = 8'h21;
  picture_data[ 4215 ] = 8'h22;
  picture_data[ 4216 ] = 8'h29;
  picture_data[ 4217 ] = 8'h62;
  picture_data[ 4218 ] = 8'h31;
  picture_data[ 4219 ] = 8'h82;
  picture_data[ 4220 ] = 8'h31;
  picture_data[ 4221 ] = 8'hC3;
  picture_data[ 4222 ] = 8'h29;
  picture_data[ 4223 ] = 8'h82;
  picture_data[ 4224 ] = 8'h31;
  picture_data[ 4225 ] = 8'hC4;
  picture_data[ 4226 ] = 8'h3A;
  picture_data[ 4227 ] = 8'h05;
  picture_data[ 4228 ] = 8'h21;
  picture_data[ 4229 ] = 8'h21;
  picture_data[ 4230 ] = 8'h39;
  picture_data[ 4231 ] = 8'hC3;
  picture_data[ 4232 ] = 8'h4A;
  picture_data[ 4233 ] = 8'h25;
  picture_data[ 4234 ] = 8'h31;
  picture_data[ 4235 ] = 8'h83;
  picture_data[ 4236 ] = 8'h31;
  picture_data[ 4237 ] = 8'h21;
  picture_data[ 4238 ] = 8'h39;
  picture_data[ 4239 ] = 8'h41;
  picture_data[ 4240 ] = 8'h41;
  picture_data[ 4241 ] = 8'hA2;
  picture_data[ 4242 ] = 8'h52;
  picture_data[ 4243 ] = 8'h03;
  picture_data[ 4244 ] = 8'hAC;
  picture_data[ 4245 ] = 8'hCE;
  picture_data[ 4246 ] = 8'hB4;
  picture_data[ 4247 ] = 8'hEF;
  picture_data[ 4248 ] = 8'hA4;
  picture_data[ 4249 ] = 8'hAF;
  picture_data[ 4250 ] = 8'hA4;
  picture_data[ 4251 ] = 8'h8F;
  picture_data[ 4252 ] = 8'h94;
  picture_data[ 4253 ] = 8'h6E;
  picture_data[ 4254 ] = 8'h8C;
  picture_data[ 4255 ] = 8'h4E;
  picture_data[ 4256 ] = 8'h5A;
  picture_data[ 4257 ] = 8'hE9;
  picture_data[ 4258 ] = 8'h73;
  picture_data[ 4259 ] = 8'hCD;
  picture_data[ 4260 ] = 8'h10;
  picture_data[ 4261 ] = 8'hE2;
  picture_data[ 4262 ] = 8'h10;
  picture_data[ 4263 ] = 8'hE3;
  picture_data[ 4264 ] = 8'h11;
  picture_data[ 4265 ] = 8'h03;
  picture_data[ 4266 ] = 8'h11;
  picture_data[ 4267 ] = 8'h03;
  picture_data[ 4268 ] = 8'h10;
  picture_data[ 4269 ] = 8'hE2;
  picture_data[ 4270 ] = 8'h19;
  picture_data[ 4271 ] = 8'h23;
  picture_data[ 4272 ] = 8'h18;
  picture_data[ 4273 ] = 8'hE3;
  picture_data[ 4274 ] = 8'h19;
  picture_data[ 4275 ] = 8'h24;
  picture_data[ 4276 ] = 8'h19;
  picture_data[ 4277 ] = 8'h03;
  picture_data[ 4278 ] = 8'h21;
  picture_data[ 4279 ] = 8'h64;
  picture_data[ 4280 ] = 8'h29;
  picture_data[ 4281 ] = 8'hA4;
  picture_data[ 4282 ] = 8'h31;
  picture_data[ 4283 ] = 8'hA5;
  picture_data[ 4284 ] = 8'h31;
  picture_data[ 4285 ] = 8'hC6;
  picture_data[ 4286 ] = 8'h31;
  picture_data[ 4287 ] = 8'hA5;
  picture_data[ 4288 ] = 8'h21;
  picture_data[ 4289 ] = 8'h43;
  picture_data[ 4290 ] = 8'h39;
  picture_data[ 4291 ] = 8'hE5;
  picture_data[ 4292 ] = 8'h21;
  picture_data[ 4293 ] = 8'h42;
  picture_data[ 4294 ] = 8'h21;
  picture_data[ 4295 ] = 8'h63;
  picture_data[ 4296 ] = 8'h21;
  picture_data[ 4297 ] = 8'h43;
  picture_data[ 4298 ] = 8'h31;
  picture_data[ 4299 ] = 8'hC5;
  picture_data[ 4300 ] = 8'h19;
  picture_data[ 4301 ] = 8'h01;
  picture_data[ 4302 ] = 8'h10;
  picture_data[ 4303 ] = 8'hC0;
  picture_data[ 4304 ] = 8'h21;
  picture_data[ 4305 ] = 8'h21;
  picture_data[ 4306 ] = 8'h29;
  picture_data[ 4307 ] = 8'h62;
  picture_data[ 4308 ] = 8'h21;
  picture_data[ 4309 ] = 8'h01;
  picture_data[ 4310 ] = 8'h21;
  picture_data[ 4311 ] = 8'h22;
  picture_data[ 4312 ] = 8'h21;
  picture_data[ 4313 ] = 8'h03;
  picture_data[ 4314 ] = 8'h29;
  picture_data[ 4315 ] = 8'h24;
  picture_data[ 4316 ] = 8'h20;
  picture_data[ 4317 ] = 8'hC2;
  picture_data[ 4318 ] = 8'h39;
  picture_data[ 4319 ] = 8'h85;
  picture_data[ 4320 ] = 8'h29;
  picture_data[ 4321 ] = 8'h03;
  picture_data[ 4322 ] = 8'h18;
  picture_data[ 4323 ] = 8'hA1;
  picture_data[ 4324 ] = 8'h20;
  picture_data[ 4325 ] = 8'hE2;
  picture_data[ 4326 ] = 8'h29;
  picture_data[ 4327 ] = 8'h02;
  picture_data[ 4328 ] = 8'h31;
  picture_data[ 4329 ] = 8'h84;
  picture_data[ 4330 ] = 8'h41;
  picture_data[ 4331 ] = 8'hE6;
  picture_data[ 4332 ] = 8'h4A;
  picture_data[ 4333 ] = 8'h27;
  picture_data[ 4334 ] = 8'h41;
  picture_data[ 4335 ] = 8'hE7;
  picture_data[ 4336 ] = 8'h39;
  picture_data[ 4337 ] = 8'hA6;
  picture_data[ 4338 ] = 8'h31;
  picture_data[ 4339 ] = 8'h85;
  picture_data[ 4340 ] = 8'h41;
  picture_data[ 4341 ] = 8'hC5;
  picture_data[ 4342 ] = 8'h31;
  picture_data[ 4343 ] = 8'h63;
  picture_data[ 4344 ] = 8'h39;
  picture_data[ 4345 ] = 8'h84;
  picture_data[ 4346 ] = 8'h41;
  picture_data[ 4347 ] = 8'hC4;
  picture_data[ 4348 ] = 8'h52;
  picture_data[ 4349 ] = 8'h88;
  picture_data[ 4350 ] = 8'h31;
  picture_data[ 4351 ] = 8'h64;
  picture_data[ 4352 ] = 8'h29;
  picture_data[ 4353 ] = 8'h64;
  picture_data[ 4354 ] = 8'h31;
  picture_data[ 4355 ] = 8'hA5;
  picture_data[ 4356 ] = 8'h29;
  picture_data[ 4357 ] = 8'h43;
  picture_data[ 4358 ] = 8'h21;
  picture_data[ 4359 ] = 8'h22;
  picture_data[ 4360 ] = 8'h21;
  picture_data[ 4361 ] = 8'h22;
  picture_data[ 4362 ] = 8'h29;
  picture_data[ 4363 ] = 8'h63;
  picture_data[ 4364 ] = 8'h31;
  picture_data[ 4365 ] = 8'hA4;
  picture_data[ 4366 ] = 8'h31;
  picture_data[ 4367 ] = 8'hC4;
  picture_data[ 4368 ] = 8'h29;
  picture_data[ 4369 ] = 8'h62;
  picture_data[ 4370 ] = 8'h31;
  picture_data[ 4371 ] = 8'hA2;
  picture_data[ 4372 ] = 8'h31;
  picture_data[ 4373 ] = 8'hA3;
  picture_data[ 4374 ] = 8'h29;
  picture_data[ 4375 ] = 8'h62;
  picture_data[ 4376 ] = 8'h29;
  picture_data[ 4377 ] = 8'h63;
  picture_data[ 4378 ] = 8'h31;
  picture_data[ 4379 ] = 8'h84;
  picture_data[ 4380 ] = 8'h21;
  picture_data[ 4381 ] = 8'h01;
  picture_data[ 4382 ] = 8'h42;
  picture_data[ 4383 ] = 8'h05;
  picture_data[ 4384 ] = 8'h29;
  picture_data[ 4385 ] = 8'h01;
  picture_data[ 4386 ] = 8'h31;
  picture_data[ 4387 ] = 8'h01;
  picture_data[ 4388 ] = 8'h51;
  picture_data[ 4389 ] = 8'h83;
  picture_data[ 4390 ] = 8'h51;
  picture_data[ 4391 ] = 8'h62;
  picture_data[ 4392 ] = 8'h51;
  picture_data[ 4393 ] = 8'hE3;
  picture_data[ 4394 ] = 8'h5A;
  picture_data[ 4395 ] = 8'h24;
  picture_data[ 4396 ] = 8'h9C;
  picture_data[ 4397 ] = 8'h4C;
  picture_data[ 4398 ] = 8'hAC;
  picture_data[ 4399 ] = 8'hEF;
  picture_data[ 4400 ] = 8'hAC;
  picture_data[ 4401 ] = 8'hF0;
  picture_data[ 4402 ] = 8'h6B;
  picture_data[ 4403 ] = 8'h29;
  picture_data[ 4404 ] = 8'h31;
  picture_data[ 4405 ] = 8'h83;
  picture_data[ 4406 ] = 8'h31;
  picture_data[ 4407 ] = 8'hC4;
  picture_data[ 4408 ] = 8'h52;
  picture_data[ 4409 ] = 8'h88;
  picture_data[ 4410 ] = 8'h42;
  picture_data[ 4411 ] = 8'h47;
  picture_data[ 4412 ] = 8'h21;
  picture_data[ 4413 ] = 8'h65;
  picture_data[ 4414 ] = 8'h10;
  picture_data[ 4415 ] = 8'hE3;
  picture_data[ 4416 ] = 8'h11;
  picture_data[ 4417 ] = 8'h03;
  picture_data[ 4418 ] = 8'h11;
  picture_data[ 4419 ] = 8'h23;
  picture_data[ 4420 ] = 8'h21;
  picture_data[ 4421 ] = 8'h64;
  picture_data[ 4422 ] = 8'h21;
  picture_data[ 4423 ] = 8'h64;
  picture_data[ 4424 ] = 8'h21;
  picture_data[ 4425 ] = 8'h85;
  picture_data[ 4426 ] = 8'h21;
  picture_data[ 4427 ] = 8'h85;
  picture_data[ 4428 ] = 8'h19;
  picture_data[ 4429 ] = 8'h23;
  picture_data[ 4430 ] = 8'h21;
  picture_data[ 4431 ] = 8'h64;
  picture_data[ 4432 ] = 8'h3A;
  picture_data[ 4433 ] = 8'h47;
  picture_data[ 4434 ] = 8'h21;
  picture_data[ 4435 ] = 8'h63;
  picture_data[ 4436 ] = 8'h18;
  picture_data[ 4437 ] = 8'hE3;
  picture_data[ 4438 ] = 8'h21;
  picture_data[ 4439 ] = 8'h23;
  picture_data[ 4440 ] = 8'h29;
  picture_data[ 4441 ] = 8'h65;
  picture_data[ 4442 ] = 8'h3A;
  picture_data[ 4443 ] = 8'h27;
  picture_data[ 4444 ] = 8'h4A;
  picture_data[ 4445 ] = 8'hC9;
  picture_data[ 4446 ] = 8'h00;
  picture_data[ 4447 ] = 8'hA0;
  picture_data[ 4448 ] = 8'h11;
  picture_data[ 4449 ] = 8'h02;
  picture_data[ 4450 ] = 8'h29;
  picture_data[ 4451 ] = 8'hA4;
  picture_data[ 4452 ] = 8'h29;
  picture_data[ 4453 ] = 8'h83;
  picture_data[ 4454 ] = 8'h31;
  picture_data[ 4455 ] = 8'hA4;
  picture_data[ 4456 ] = 8'h29;
  picture_data[ 4457 ] = 8'h42;
  picture_data[ 4458 ] = 8'h31;
  picture_data[ 4459 ] = 8'hA3;
  picture_data[ 4460 ] = 8'h29;
  picture_data[ 4461 ] = 8'h22;
  picture_data[ 4462 ] = 8'h29;
  picture_data[ 4463 ] = 8'h43;
  picture_data[ 4464 ] = 8'h18;
  picture_data[ 4465 ] = 8'hC1;
  picture_data[ 4466 ] = 8'h21;
  picture_data[ 4467 ] = 8'h03;
  picture_data[ 4468 ] = 8'h31;
  picture_data[ 4469 ] = 8'h43;
  picture_data[ 4470 ] = 8'h10;
  picture_data[ 4471 ] = 8'h60;
  picture_data[ 4472 ] = 8'h29;
  picture_data[ 4473 ] = 8'h23;
  picture_data[ 4474 ] = 8'h41;
  picture_data[ 4475 ] = 8'hC5;
  picture_data[ 4476 ] = 8'h31;
  picture_data[ 4477 ] = 8'h64;
  picture_data[ 4478 ] = 8'h39;
  picture_data[ 4479 ] = 8'hA4;
  picture_data[ 4480 ] = 8'h52;
  picture_data[ 4481 ] = 8'h47;
  picture_data[ 4482 ] = 8'h5A;
  picture_data[ 4483 ] = 8'hA9;
  picture_data[ 4484 ] = 8'h31;
  picture_data[ 4485 ] = 8'h84;
  picture_data[ 4486 ] = 8'h39;
  picture_data[ 4487 ] = 8'hA5;
  picture_data[ 4488 ] = 8'h31;
  picture_data[ 4489 ] = 8'h84;
  picture_data[ 4490 ] = 8'h41;
  picture_data[ 4491 ] = 8'hE6;
  picture_data[ 4492 ] = 8'h39;
  picture_data[ 4493 ] = 8'h84;
  picture_data[ 4494 ] = 8'h39;
  picture_data[ 4495 ] = 8'h83;
  picture_data[ 4496 ] = 8'h39;
  picture_data[ 4497 ] = 8'hA3;
  picture_data[ 4498 ] = 8'h41;
  picture_data[ 4499 ] = 8'hE5;
  picture_data[ 4500 ] = 8'h42;
  picture_data[ 4501 ] = 8'h05;
  picture_data[ 4502 ] = 8'h31;
  picture_data[ 4503 ] = 8'h84;
  picture_data[ 4504 ] = 8'h29;
  picture_data[ 4505 ] = 8'h64;
  picture_data[ 4506 ] = 8'h29;
  picture_data[ 4507 ] = 8'h84;
  picture_data[ 4508 ] = 8'h29;
  picture_data[ 4509 ] = 8'h43;
  picture_data[ 4510 ] = 8'h21;
  picture_data[ 4511 ] = 8'h22;
  picture_data[ 4512 ] = 8'h19;
  picture_data[ 4513 ] = 8'h02;
  picture_data[ 4514 ] = 8'h21;
  picture_data[ 4515 ] = 8'h02;
  picture_data[ 4516 ] = 8'h29;
  picture_data[ 4517 ] = 8'h63;
  picture_data[ 4518 ] = 8'h31;
  picture_data[ 4519 ] = 8'hC4;
  picture_data[ 4520 ] = 8'h31;
  picture_data[ 4521 ] = 8'h83;
  picture_data[ 4522 ] = 8'h39;
  picture_data[ 4523 ] = 8'hE4;
  picture_data[ 4524 ] = 8'h39;
  picture_data[ 4525 ] = 8'hE4;
  picture_data[ 4526 ] = 8'h42;
  picture_data[ 4527 ] = 8'h05;
  picture_data[ 4528 ] = 8'h31;
  picture_data[ 4529 ] = 8'h84;
  picture_data[ 4530 ] = 8'h21;
  picture_data[ 4531 ] = 8'h02;
  picture_data[ 4532 ] = 8'h20;
  picture_data[ 4533 ] = 8'hE1;
  picture_data[ 4534 ] = 8'h29;
  picture_data[ 4535 ] = 8'h22;
  picture_data[ 4536 ] = 8'h20;
  picture_data[ 4537 ] = 8'hC0;
  picture_data[ 4538 ] = 8'h41;
  picture_data[ 4539 ] = 8'h21;
  picture_data[ 4540 ] = 8'h59;
  picture_data[ 4541 ] = 8'h63;
  picture_data[ 4542 ] = 8'h69;
  picture_data[ 4543 ] = 8'hC4;
  picture_data[ 4544 ] = 8'h72;
  picture_data[ 4545 ] = 8'h65;
  picture_data[ 4546 ] = 8'h5A;
  picture_data[ 4547 ] = 8'h03;
  picture_data[ 4548 ] = 8'h8B;
  picture_data[ 4549 ] = 8'hAA;
  picture_data[ 4550 ] = 8'hB5;
  picture_data[ 4551 ] = 8'h30;
  picture_data[ 4552 ] = 8'h94;
  picture_data[ 4553 ] = 8'h2D;
  picture_data[ 4554 ] = 8'h5A;
  picture_data[ 4555 ] = 8'h87;
  picture_data[ 4556 ] = 8'h4A;
  picture_data[ 4557 ] = 8'h47;
  picture_data[ 4558 ] = 8'h52;
  picture_data[ 4559 ] = 8'hE9;
  picture_data[ 4560 ] = 8'h21;
  picture_data[ 4561 ] = 8'h03;
  picture_data[ 4562 ] = 8'h10;
  picture_data[ 4563 ] = 8'h61;
  picture_data[ 4564 ] = 8'h21;
  picture_data[ 4565 ] = 8'h45;
  picture_data[ 4566 ] = 8'h19;
  picture_data[ 4567 ] = 8'h25;
  picture_data[ 4568 ] = 8'h21;
  picture_data[ 4569 ] = 8'h65;
  picture_data[ 4570 ] = 8'h21;
  picture_data[ 4571 ] = 8'h85;
  picture_data[ 4572 ] = 8'h29;
  picture_data[ 4573 ] = 8'hA4;
  picture_data[ 4574 ] = 8'h11;
  picture_data[ 4575 ] = 8'h02;
  picture_data[ 4576 ] = 8'h19;
  picture_data[ 4577 ] = 8'h23;
  picture_data[ 4578 ] = 8'h29;
  picture_data[ 4579 ] = 8'hA5;
  picture_data[ 4580 ] = 8'h19;
  picture_data[ 4581 ] = 8'h44;
  picture_data[ 4582 ] = 8'h21;
  picture_data[ 4583 ] = 8'h64;
  picture_data[ 4584 ] = 8'h11;
  picture_data[ 4585 ] = 8'h22;
  picture_data[ 4586 ] = 8'h29;
  picture_data[ 4587 ] = 8'hC5;
  picture_data[ 4588 ] = 8'h29;
  picture_data[ 4589 ] = 8'hA5;
  picture_data[ 4590 ] = 8'h21;
  picture_data[ 4591 ] = 8'h24;
  picture_data[ 4592 ] = 8'h21;
  picture_data[ 4593 ] = 8'h85;
  picture_data[ 4594 ] = 8'h29;
  picture_data[ 4595 ] = 8'hC6;
  picture_data[ 4596 ] = 8'h19;
  picture_data[ 4597 ] = 8'h84;
  picture_data[ 4598 ] = 8'h09;
  picture_data[ 4599 ] = 8'h02;
  picture_data[ 4600 ] = 8'h00;
  picture_data[ 4601 ] = 8'hA0;
  picture_data[ 4602 ] = 8'h21;
  picture_data[ 4603 ] = 8'h84;
  picture_data[ 4604 ] = 8'h21;
  picture_data[ 4605 ] = 8'h42;
  picture_data[ 4606 ] = 8'h21;
  picture_data[ 4607 ] = 8'h02;
  picture_data[ 4608 ] = 8'h29;
  picture_data[ 4609 ] = 8'h02;
  picture_data[ 4610 ] = 8'h31;
  picture_data[ 4611 ] = 8'h23;
  picture_data[ 4612 ] = 8'h18;
  picture_data[ 4613 ] = 8'hC1;
  picture_data[ 4614 ] = 8'h20;
  picture_data[ 4615 ] = 8'hE2;
  picture_data[ 4616 ] = 8'h29;
  picture_data[ 4617 ] = 8'h43;
  picture_data[ 4618 ] = 8'h21;
  picture_data[ 4619 ] = 8'h22;
  picture_data[ 4620 ] = 8'h29;
  picture_data[ 4621 ] = 8'h43;
  picture_data[ 4622 ] = 8'h31;
  picture_data[ 4623 ] = 8'h63;
  picture_data[ 4624 ] = 8'h20;
  picture_data[ 4625 ] = 8'hE2;
  picture_data[ 4626 ] = 8'h31;
  picture_data[ 4627 ] = 8'h44;
  picture_data[ 4628 ] = 8'h31;
  picture_data[ 4629 ] = 8'h63;
  picture_data[ 4630 ] = 8'h29;
  picture_data[ 4631 ] = 8'h02;
  picture_data[ 4632 ] = 8'h4A;
  picture_data[ 4633 ] = 8'h06;
  picture_data[ 4634 ] = 8'h4A;
  picture_data[ 4635 ] = 8'h27;
  picture_data[ 4636 ] = 8'h31;
  picture_data[ 4637 ] = 8'h84;
  picture_data[ 4638 ] = 8'h39;
  picture_data[ 4639 ] = 8'hA5;
  picture_data[ 4640 ] = 8'h39;
  picture_data[ 4641 ] = 8'hC5;
  picture_data[ 4642 ] = 8'h41;
  picture_data[ 4643 ] = 8'hE6;
  picture_data[ 4644 ] = 8'h39;
  picture_data[ 4645 ] = 8'hA4;
  picture_data[ 4646 ] = 8'h39;
  picture_data[ 4647 ] = 8'hE4;
  picture_data[ 4648 ] = 8'h31;
  picture_data[ 4649 ] = 8'h62;
  picture_data[ 4650 ] = 8'h39;
  picture_data[ 4651 ] = 8'hC4;
  picture_data[ 4652 ] = 8'h31;
  picture_data[ 4653 ] = 8'h83;
  picture_data[ 4654 ] = 8'h31;
  picture_data[ 4655 ] = 8'h64;
  picture_data[ 4656 ] = 8'h21;
  picture_data[ 4657 ] = 8'h02;
  picture_data[ 4658 ] = 8'h18;
  picture_data[ 4659 ] = 8'hC1;
  picture_data[ 4660 ] = 8'h19;
  picture_data[ 4661 ] = 8'h01;
  picture_data[ 4662 ] = 8'h29;
  picture_data[ 4663 ] = 8'h62;
  picture_data[ 4664 ] = 8'h29;
  picture_data[ 4665 ] = 8'h63;
  picture_data[ 4666 ] = 8'h21;
  picture_data[ 4667 ] = 8'h23;
  picture_data[ 4668 ] = 8'h21;
  picture_data[ 4669 ] = 8'h23;
  picture_data[ 4670 ] = 8'h29;
  picture_data[ 4671 ] = 8'h63;
  picture_data[ 4672 ] = 8'h31;
  picture_data[ 4673 ] = 8'hA3;
  picture_data[ 4674 ] = 8'h39;
  picture_data[ 4675 ] = 8'hE4;
  picture_data[ 4676 ] = 8'h39;
  picture_data[ 4677 ] = 8'hE4;
  picture_data[ 4678 ] = 8'h42;
  picture_data[ 4679 ] = 8'h05;
  picture_data[ 4680 ] = 8'h31;
  picture_data[ 4681 ] = 8'h84;
  picture_data[ 4682 ] = 8'h18;
  picture_data[ 4683 ] = 8'hC2;
  picture_data[ 4684 ] = 8'h20;
  picture_data[ 4685 ] = 8'hE2;
  picture_data[ 4686 ] = 8'h18;
  picture_data[ 4687 ] = 8'hA0;
  picture_data[ 4688 ] = 8'h20;
  picture_data[ 4689 ] = 8'hC0;
  picture_data[ 4690 ] = 8'h51;
  picture_data[ 4691 ] = 8'hA4;
  picture_data[ 4692 ] = 8'h71;
  picture_data[ 4693 ] = 8'hA5;
  picture_data[ 4694 ] = 8'h79;
  picture_data[ 4695 ] = 8'hE5;
  picture_data[ 4696 ] = 8'h72;
  picture_data[ 4697 ] = 8'h04;
  picture_data[ 4698 ] = 8'h6A;
  picture_data[ 4699 ] = 8'h24;
  picture_data[ 4700 ] = 8'h59;
  picture_data[ 4701 ] = 8'hE3;
  picture_data[ 4702 ] = 8'h41;
  picture_data[ 4703 ] = 8'h41;
  picture_data[ 4704 ] = 8'h5A;
  picture_data[ 4705 ] = 8'h25;
  picture_data[ 4706 ] = 8'h93;
  picture_data[ 4707 ] = 8'hED;
  picture_data[ 4708 ] = 8'h5A;
  picture_data[ 4709 ] = 8'h88;
  picture_data[ 4710 ] = 8'h39;
  picture_data[ 4711 ] = 8'hA4;
  picture_data[ 4712 ] = 8'h18;
  picture_data[ 4713 ] = 8'h82;
  picture_data[ 4714 ] = 8'h29;
  picture_data[ 4715 ] = 8'h65;
  picture_data[ 4716 ] = 8'h21;
  picture_data[ 4717 ] = 8'h46;
  picture_data[ 4718 ] = 8'h21;
  picture_data[ 4719 ] = 8'h46;
  picture_data[ 4720 ] = 8'h19;
  picture_data[ 4721 ] = 8'h24;
  picture_data[ 4722 ] = 8'h08;
  picture_data[ 4723 ] = 8'hE2;
  picture_data[ 4724 ] = 8'h00;
  picture_data[ 4725 ] = 8'h80;
  picture_data[ 4726 ] = 8'h08;
  picture_data[ 4727 ] = 8'hA1;
  picture_data[ 4728 ] = 8'h08;
  picture_data[ 4729 ] = 8'hA1;
  picture_data[ 4730 ] = 8'h19;
  picture_data[ 4731 ] = 8'h23;
  picture_data[ 4732 ] = 8'h19;
  picture_data[ 4733 ] = 8'h44;
  picture_data[ 4734 ] = 8'h19;
  picture_data[ 4735 ] = 8'h23;
  picture_data[ 4736 ] = 8'h21;
  picture_data[ 4737 ] = 8'h85;
  picture_data[ 4738 ] = 8'h21;
  picture_data[ 4739 ] = 8'h84;
  picture_data[ 4740 ] = 8'h21;
  picture_data[ 4741 ] = 8'h85;
  picture_data[ 4742 ] = 8'h11;
  picture_data[ 4743 ] = 8'h03;
  picture_data[ 4744 ] = 8'h11;
  picture_data[ 4745 ] = 8'h03;
  picture_data[ 4746 ] = 8'h11;
  picture_data[ 4747 ] = 8'h23;
  picture_data[ 4748 ] = 8'h32;
  picture_data[ 4749 ] = 8'h48;
  picture_data[ 4750 ] = 8'h21;
  picture_data[ 4751 ] = 8'hC5;
  picture_data[ 4752 ] = 8'h09;
  picture_data[ 4753 ] = 8'h02;
  picture_data[ 4754 ] = 8'h11;
  picture_data[ 4755 ] = 8'h22;
  picture_data[ 4756 ] = 8'h21;
  picture_data[ 4757 ] = 8'h43;
  picture_data[ 4758 ] = 8'h21;
  picture_data[ 4759 ] = 8'h22;
  picture_data[ 4760 ] = 8'h29;
  picture_data[ 4761 ] = 8'h43;
  picture_data[ 4762 ] = 8'h20;
  picture_data[ 4763 ] = 8'hE2;
  picture_data[ 4764 ] = 8'h21;
  picture_data[ 4765 ] = 8'h03;
  picture_data[ 4766 ] = 8'h20;
  picture_data[ 4767 ] = 8'hE2;
  picture_data[ 4768 ] = 8'h31;
  picture_data[ 4769 ] = 8'h83;
  picture_data[ 4770 ] = 8'h31;
  picture_data[ 4771 ] = 8'h83;
  picture_data[ 4772 ] = 8'h21;
  picture_data[ 4773 ] = 8'h02;
  picture_data[ 4774 ] = 8'h31;
  picture_data[ 4775 ] = 8'h84;
  picture_data[ 4776 ] = 8'h39;
  picture_data[ 4777 ] = 8'hA5;
  picture_data[ 4778 ] = 8'h20;
  picture_data[ 4779 ] = 8'hE2;
  picture_data[ 4780 ] = 8'h21;
  picture_data[ 4781 ] = 8'h02;
  picture_data[ 4782 ] = 8'h31;
  picture_data[ 4783 ] = 8'h64;
  picture_data[ 4784 ] = 8'h39;
  picture_data[ 4785 ] = 8'h84;
  picture_data[ 4786 ] = 8'h4A;
  picture_data[ 4787 ] = 8'h06;
  picture_data[ 4788 ] = 8'h42;
  picture_data[ 4789 ] = 8'h06;
  picture_data[ 4790 ] = 8'h42;
  picture_data[ 4791 ] = 8'h06;
  picture_data[ 4792 ] = 8'h39;
  picture_data[ 4793 ] = 8'hC5;
  picture_data[ 4794 ] = 8'h31;
  picture_data[ 4795 ] = 8'hA4;
  picture_data[ 4796 ] = 8'h42;
  picture_data[ 4797 ] = 8'h05;
  picture_data[ 4798 ] = 8'h29;
  picture_data[ 4799 ] = 8'h42;
  picture_data[ 4800 ] = 8'h31;
  picture_data[ 4801 ] = 8'hA4;
  picture_data[ 4802 ] = 8'h31;
  picture_data[ 4803 ] = 8'h63;
  picture_data[ 4804 ] = 8'h31;
  picture_data[ 4805 ] = 8'h83;
  picture_data[ 4806 ] = 8'h31;
  picture_data[ 4807 ] = 8'h84;
  picture_data[ 4808 ] = 8'h29;
  picture_data[ 4809 ] = 8'h63;
  picture_data[ 4810 ] = 8'h21;
  picture_data[ 4811 ] = 8'h22;
  picture_data[ 4812 ] = 8'h21;
  picture_data[ 4813 ] = 8'h42;
  picture_data[ 4814 ] = 8'h29;
  picture_data[ 4815 ] = 8'h83;
  picture_data[ 4816 ] = 8'h31;
  picture_data[ 4817 ] = 8'hA4;
  picture_data[ 4818 ] = 8'h31;
  picture_data[ 4819 ] = 8'hA4;
  picture_data[ 4820 ] = 8'h29;
  picture_data[ 4821 ] = 8'h63;
  picture_data[ 4822 ] = 8'h21;
  picture_data[ 4823 ] = 8'h42;
  picture_data[ 4824 ] = 8'h21;
  picture_data[ 4825 ] = 8'h42;
  picture_data[ 4826 ] = 8'h29;
  picture_data[ 4827 ] = 8'h62;
  picture_data[ 4828 ] = 8'h21;
  picture_data[ 4829 ] = 8'h21;
  picture_data[ 4830 ] = 8'h18;
  picture_data[ 4831 ] = 8'hE1;
  picture_data[ 4832 ] = 8'h21;
  picture_data[ 4833 ] = 8'h02;
  picture_data[ 4834 ] = 8'h18;
  picture_data[ 4835 ] = 8'hC1;
  picture_data[ 4836 ] = 8'h20;
  picture_data[ 4837 ] = 8'hC1;
  picture_data[ 4838 ] = 8'h20;
  picture_data[ 4839 ] = 8'hE1;
  picture_data[ 4840 ] = 8'h31;
  picture_data[ 4841 ] = 8'h43;
  picture_data[ 4842 ] = 8'h30;
  picture_data[ 4843 ] = 8'hE1;
  picture_data[ 4844 ] = 8'h69;
  picture_data[ 4845 ] = 8'hC5;
  picture_data[ 4846 ] = 8'h8A;
  picture_data[ 4847 ] = 8'h87;
  picture_data[ 4848 ] = 8'h6A;
  picture_data[ 4849 ] = 8'h04;
  picture_data[ 4850 ] = 8'h72;
  picture_data[ 4851 ] = 8'hA6;
  picture_data[ 4852 ] = 8'h51;
  picture_data[ 4853 ] = 8'hA2;
  picture_data[ 4854 ] = 8'h51;
  picture_data[ 4855 ] = 8'h82;
  picture_data[ 4856 ] = 8'h59;
  picture_data[ 4857 ] = 8'hE4;
  picture_data[ 4858 ] = 8'h6A;
  picture_data[ 4859 ] = 8'h67;
  picture_data[ 4860 ] = 8'h49;
  picture_data[ 4861 ] = 8'hC4;
  picture_data[ 4862 ] = 8'h52;
  picture_data[ 4863 ] = 8'h26;
  picture_data[ 4864 ] = 8'h29;
  picture_data[ 4865 ] = 8'h66;
  picture_data[ 4866 ] = 8'h19;
  picture_data[ 4867 ] = 8'h04;
  picture_data[ 4868 ] = 8'h00;
  picture_data[ 4869 ] = 8'h41;
  picture_data[ 4870 ] = 8'h00;
  picture_data[ 4871 ] = 8'h41;
  picture_data[ 4872 ] = 8'h00;
  picture_data[ 4873 ] = 8'hA2;
  picture_data[ 4874 ] = 8'h11;
  picture_data[ 4875 ] = 8'h04;
  picture_data[ 4876 ] = 8'h11;
  picture_data[ 4877 ] = 8'h04;
  picture_data[ 4878 ] = 8'h19;
  picture_data[ 4879 ] = 8'h24;
  picture_data[ 4880 ] = 8'h19;
  picture_data[ 4881 ] = 8'h03;
  picture_data[ 4882 ] = 8'h19;
  picture_data[ 4883 ] = 8'h03;
  picture_data[ 4884 ] = 8'h21;
  picture_data[ 4885 ] = 8'h44;
  picture_data[ 4886 ] = 8'h29;
  picture_data[ 4887 ] = 8'h86;
  picture_data[ 4888 ] = 8'h19;
  picture_data[ 4889 ] = 8'h24;
  picture_data[ 4890 ] = 8'h21;
  picture_data[ 4891 ] = 8'h44;
  picture_data[ 4892 ] = 8'h19;
  picture_data[ 4893 ] = 8'h03;
  picture_data[ 4894 ] = 8'h11;
  picture_data[ 4895 ] = 8'h02;
  picture_data[ 4896 ] = 8'h00;
  picture_data[ 4897 ] = 8'hE2;
  picture_data[ 4898 ] = 8'h19;
  picture_data[ 4899 ] = 8'hE6;
  picture_data[ 4900 ] = 8'h6C;
  picture_data[ 4901 ] = 8'h2F;
  picture_data[ 4902 ] = 8'h32;
  picture_data[ 4903 ] = 8'h67;
  picture_data[ 4904 ] = 8'h19;
  picture_data[ 4905 ] = 8'h64;
  picture_data[ 4906 ] = 8'h21;
  picture_data[ 4907 ] = 8'h84;
  picture_data[ 4908 ] = 8'h10;
  picture_data[ 4909 ] = 8'hE2;
  picture_data[ 4910 ] = 8'h31;
  picture_data[ 4911 ] = 8'hC5;
  picture_data[ 4912 ] = 8'h31;
  picture_data[ 4913 ] = 8'h85;
  picture_data[ 4914 ] = 8'h18;
  picture_data[ 4915 ] = 8'hE2;
  picture_data[ 4916 ] = 8'h20;
  picture_data[ 4917 ] = 8'hE2;
  picture_data[ 4918 ] = 8'h21;
  picture_data[ 4919 ] = 8'h02;
  picture_data[ 4920 ] = 8'h21;
  picture_data[ 4921 ] = 8'h02;
  picture_data[ 4922 ] = 8'h21;
  picture_data[ 4923 ] = 8'h02;
  picture_data[ 4924 ] = 8'h29;
  picture_data[ 4925 ] = 8'h64;
  picture_data[ 4926 ] = 8'h29;
  picture_data[ 4927 ] = 8'h43;
  picture_data[ 4928 ] = 8'h42;
  picture_data[ 4929 ] = 8'h06;
  picture_data[ 4930 ] = 8'h4A;
  picture_data[ 4931 ] = 8'h26;
  picture_data[ 4932 ] = 8'h31;
  picture_data[ 4933 ] = 8'h64;
  picture_data[ 4934 ] = 8'h31;
  picture_data[ 4935 ] = 8'h85;
  picture_data[ 4936 ] = 8'h29;
  picture_data[ 4937 ] = 8'h44;
  picture_data[ 4938 ] = 8'h41;
  picture_data[ 4939 ] = 8'hE6;
  picture_data[ 4940 ] = 8'h4A;
  picture_data[ 4941 ] = 8'h27;
  picture_data[ 4942 ] = 8'h52;
  picture_data[ 4943 ] = 8'h88;
  picture_data[ 4944 ] = 8'h41;
  picture_data[ 4945 ] = 8'hE5;
  picture_data[ 4946 ] = 8'h21;
  picture_data[ 4947 ] = 8'h21;
  picture_data[ 4948 ] = 8'h29;
  picture_data[ 4949 ] = 8'h42;
  picture_data[ 4950 ] = 8'h29;
  picture_data[ 4951 ] = 8'h62;
  picture_data[ 4952 ] = 8'h39;
  picture_data[ 4953 ] = 8'hC4;
  picture_data[ 4954 ] = 8'h29;
  picture_data[ 4955 ] = 8'h43;
  picture_data[ 4956 ] = 8'h21;
  picture_data[ 4957 ] = 8'h22;
  picture_data[ 4958 ] = 8'h29;
  picture_data[ 4959 ] = 8'h43;
  picture_data[ 4960 ] = 8'h29;
  picture_data[ 4961 ] = 8'h83;
  picture_data[ 4962 ] = 8'h21;
  picture_data[ 4963 ] = 8'h43;
  picture_data[ 4964 ] = 8'h29;
  picture_data[ 4965 ] = 8'h63;
  picture_data[ 4966 ] = 8'h31;
  picture_data[ 4967 ] = 8'hE5;
  picture_data[ 4968 ] = 8'h29;
  picture_data[ 4969 ] = 8'hA4;
  picture_data[ 4970 ] = 8'h21;
  picture_data[ 4971 ] = 8'h42;
  picture_data[ 4972 ] = 8'h21;
  picture_data[ 4973 ] = 8'h42;
  picture_data[ 4974 ] = 8'h39;
  picture_data[ 4975 ] = 8'hE5;
  picture_data[ 4976 ] = 8'h39;
  picture_data[ 4977 ] = 8'hE4;
  picture_data[ 4978 ] = 8'h29;
  picture_data[ 4979 ] = 8'h83;
  picture_data[ 4980 ] = 8'h39;
  picture_data[ 4981 ] = 8'hC4;
  picture_data[ 4982 ] = 8'h18;
  picture_data[ 4983 ] = 8'hE1;
  picture_data[ 4984 ] = 8'h41;
  picture_data[ 4985 ] = 8'hE5;
  picture_data[ 4986 ] = 8'h39;
  picture_data[ 4987 ] = 8'hA4;
  picture_data[ 4988 ] = 8'h29;
  picture_data[ 4989 ] = 8'h22;
  picture_data[ 4990 ] = 8'h29;
  picture_data[ 4991 ] = 8'h22;
  picture_data[ 4992 ] = 8'h31;
  picture_data[ 4993 ] = 8'h63;
  picture_data[ 4994 ] = 8'h39;
  picture_data[ 4995 ] = 8'h63;
  picture_data[ 4996 ] = 8'h49;
  picture_data[ 4997 ] = 8'h83;
  picture_data[ 4998 ] = 8'h62;
  picture_data[ 4999 ] = 8'h45;
  picture_data[ 5000 ] = 8'h62;
  picture_data[ 5001 ] = 8'h65;
  picture_data[ 5002 ] = 8'h6A;
  picture_data[ 5003 ] = 8'h85;
  picture_data[ 5004 ] = 8'h6A;
  picture_data[ 5005 ] = 8'h85;
  picture_data[ 5006 ] = 8'h62;
  picture_data[ 5007 ] = 8'h44;
  picture_data[ 5008 ] = 8'h5A;
  picture_data[ 5009 ] = 8'h04;
  picture_data[ 5010 ] = 8'h6A;
  picture_data[ 5011 ] = 8'h66;
  picture_data[ 5012 ] = 8'h62;
  picture_data[ 5013 ] = 8'h46;
  picture_data[ 5014 ] = 8'h6A;
  picture_data[ 5015 ] = 8'h46;
  picture_data[ 5016 ] = 8'h10;
  picture_data[ 5017 ] = 8'hA4;
  picture_data[ 5018 ] = 8'h10;
  picture_data[ 5019 ] = 8'hC4;
  picture_data[ 5020 ] = 8'h08;
  picture_data[ 5021 ] = 8'h83;
  picture_data[ 5022 ] = 8'h08;
  picture_data[ 5023 ] = 8'hC3;
  picture_data[ 5024 ] = 8'h19;
  picture_data[ 5025 ] = 8'h45;
  picture_data[ 5026 ] = 8'h11;
  picture_data[ 5027 ] = 8'h25;
  picture_data[ 5028 ] = 8'h08;
  picture_data[ 5029 ] = 8'h83;
  picture_data[ 5030 ] = 8'h00;
  picture_data[ 5031 ] = 8'h42;
  picture_data[ 5032 ] = 8'h10;
  picture_data[ 5033 ] = 8'hC2;
  picture_data[ 5034 ] = 8'h08;
  picture_data[ 5035 ] = 8'h81;
  picture_data[ 5036 ] = 8'h21;
  picture_data[ 5037 ] = 8'h24;
  picture_data[ 5038 ] = 8'h18;
  picture_data[ 5039 ] = 8'hE4;
  picture_data[ 5040 ] = 8'h21;
  picture_data[ 5041 ] = 8'h45;
  picture_data[ 5042 ] = 8'h21;
  picture_data[ 5043 ] = 8'h65;
  picture_data[ 5044 ] = 8'h19;
  picture_data[ 5045 ] = 8'h23;
  picture_data[ 5046 ] = 8'h29;
  picture_data[ 5047 ] = 8'hC6;
  picture_data[ 5048 ] = 8'h01;
  picture_data[ 5049 ] = 8'h02;
  picture_data[ 5050 ] = 8'h19;
  picture_data[ 5051 ] = 8'hC6;
  picture_data[ 5052 ] = 8'h2A;
  picture_data[ 5053 ] = 8'h47;
  picture_data[ 5054 ] = 8'h11;
  picture_data[ 5055 ] = 8'h64;
  picture_data[ 5056 ] = 8'h32;
  picture_data[ 5057 ] = 8'h27;
  picture_data[ 5058 ] = 8'h08;
  picture_data[ 5059 ] = 8'hE2;
  picture_data[ 5060 ] = 8'h10;
  picture_data[ 5061 ] = 8'hE2;
  picture_data[ 5062 ] = 8'h21;
  picture_data[ 5063 ] = 8'h43;
  picture_data[ 5064 ] = 8'h21;
  picture_data[ 5065 ] = 8'h23;
  picture_data[ 5066 ] = 8'h18;
  picture_data[ 5067 ] = 8'hE2;
  picture_data[ 5068 ] = 8'h18;
  picture_data[ 5069 ] = 8'hE2;
  picture_data[ 5070 ] = 8'h18;
  picture_data[ 5071 ] = 8'hE2;
  picture_data[ 5072 ] = 8'h21;
  picture_data[ 5073 ] = 8'h22;
  picture_data[ 5074 ] = 8'h18;
  picture_data[ 5075 ] = 8'hE1;
  picture_data[ 5076 ] = 8'h18;
  picture_data[ 5077 ] = 8'hE2;
  picture_data[ 5078 ] = 8'h21;
  picture_data[ 5079 ] = 8'h23;
  picture_data[ 5080 ] = 8'h21;
  picture_data[ 5081 ] = 8'h22;
  picture_data[ 5082 ] = 8'h39;
  picture_data[ 5083 ] = 8'hC4;
  picture_data[ 5084 ] = 8'h31;
  picture_data[ 5085 ] = 8'h84;
  picture_data[ 5086 ] = 8'h20;
  picture_data[ 5087 ] = 8'hC2;
  picture_data[ 5088 ] = 8'h31;
  picture_data[ 5089 ] = 8'h44;
  picture_data[ 5090 ] = 8'h29;
  picture_data[ 5091 ] = 8'h02;
  picture_data[ 5092 ] = 8'h39;
  picture_data[ 5093 ] = 8'hA4;
  picture_data[ 5094 ] = 8'h4A;
  picture_data[ 5095 ] = 8'h25;
  picture_data[ 5096 ] = 8'h31;
  picture_data[ 5097 ] = 8'h61;
  picture_data[ 5098 ] = 8'h41;
  picture_data[ 5099 ] = 8'hE3;
  picture_data[ 5100 ] = 8'h29;
  picture_data[ 5101 ] = 8'h21;
  picture_data[ 5102 ] = 8'h31;
  picture_data[ 5103 ] = 8'h62;
  picture_data[ 5104 ] = 8'h31;
  picture_data[ 5105 ] = 8'hC4;
  picture_data[ 5106 ] = 8'h31;
  picture_data[ 5107 ] = 8'hC4;
  picture_data[ 5108 ] = 8'h29;
  picture_data[ 5109 ] = 8'h83;
  picture_data[ 5110 ] = 8'h21;
  picture_data[ 5111 ] = 8'h42;
  picture_data[ 5112 ] = 8'h21;
  picture_data[ 5113 ] = 8'h22;
  picture_data[ 5114 ] = 8'h29;
  picture_data[ 5115 ] = 8'h83;
  picture_data[ 5116 ] = 8'h31;
  picture_data[ 5117 ] = 8'hA4;
  picture_data[ 5118 ] = 8'h29;
  picture_data[ 5119 ] = 8'h83;
  picture_data[ 5120 ] = 8'h31;
  picture_data[ 5121 ] = 8'hE4;
  picture_data[ 5122 ] = 8'h3A;
  picture_data[ 5123 ] = 8'h05;
  picture_data[ 5124 ] = 8'h31;
  picture_data[ 5125 ] = 8'hA3;
  picture_data[ 5126 ] = 8'h3A;
  picture_data[ 5127 ] = 8'h05;
  picture_data[ 5128 ] = 8'h3A;
  picture_data[ 5129 ] = 8'h05;
  picture_data[ 5130 ] = 8'h39;
  picture_data[ 5131 ] = 8'hC4;
  picture_data[ 5132 ] = 8'h39;
  picture_data[ 5133 ] = 8'hC4;
  picture_data[ 5134 ] = 8'h39;
  picture_data[ 5135 ] = 8'hC4;
  picture_data[ 5136 ] = 8'h39;
  picture_data[ 5137 ] = 8'hC4;
  picture_data[ 5138 ] = 8'h39;
  picture_data[ 5139 ] = 8'hA4;
  picture_data[ 5140 ] = 8'h31;
  picture_data[ 5141 ] = 8'h83;
  picture_data[ 5142 ] = 8'h31;
  picture_data[ 5143 ] = 8'h62;
  picture_data[ 5144 ] = 8'h31;
  picture_data[ 5145 ] = 8'h63;
  picture_data[ 5146 ] = 8'h41;
  picture_data[ 5147 ] = 8'hC4;
  picture_data[ 5148 ] = 8'h41;
  picture_data[ 5149 ] = 8'hE4;
  picture_data[ 5150 ] = 8'h39;
  picture_data[ 5151 ] = 8'h61;
  picture_data[ 5152 ] = 8'h41;
  picture_data[ 5153 ] = 8'hC2;
  picture_data[ 5154 ] = 8'h5A;
  picture_data[ 5155 ] = 8'h44;
  picture_data[ 5156 ] = 8'h62;
  picture_data[ 5157 ] = 8'h64;
  picture_data[ 5158 ] = 8'h49;
  picture_data[ 5159 ] = 8'h81;
  picture_data[ 5160 ] = 8'h51;
  picture_data[ 5161 ] = 8'hC3;
  picture_data[ 5162 ] = 8'h5A;
  picture_data[ 5163 ] = 8'h04;
  picture_data[ 5164 ] = 8'h59;
  picture_data[ 5165 ] = 8'hC4;
  picture_data[ 5166 ] = 8'h62;
  picture_data[ 5167 ] = 8'h25;
  picture_data[ 5168 ] = 8'h10;
  picture_data[ 5169 ] = 8'hC5;
  picture_data[ 5170 ] = 8'h08;
  picture_data[ 5171 ] = 8'hA4;
  picture_data[ 5172 ] = 8'h21;
  picture_data[ 5173 ] = 8'h46;
  picture_data[ 5174 ] = 8'h29;
  picture_data[ 5175 ] = 8'h87;
  picture_data[ 5176 ] = 8'h08;
  picture_data[ 5177 ] = 8'hA3;
  picture_data[ 5178 ] = 8'h00;
  picture_data[ 5179 ] = 8'h62;
  picture_data[ 5180 ] = 8'h10;
  picture_data[ 5181 ] = 8'hC5;
  picture_data[ 5182 ] = 8'h08;
  picture_data[ 5183 ] = 8'hA4;
  picture_data[ 5184 ] = 8'h19;
  picture_data[ 5185 ] = 8'h25;
  picture_data[ 5186 ] = 8'h19;
  picture_data[ 5187 ] = 8'h03;
  picture_data[ 5188 ] = 8'h10;
  picture_data[ 5189 ] = 8'hA2;
  picture_data[ 5190 ] = 8'h10;
  picture_data[ 5191 ] = 8'hC3;
  picture_data[ 5192 ] = 8'h19;
  picture_data[ 5193 ] = 8'h03;
  picture_data[ 5194 ] = 8'h29;
  picture_data[ 5195 ] = 8'h65;
  picture_data[ 5196 ] = 8'h19;
  picture_data[ 5197 ] = 8'h03;
  picture_data[ 5198 ] = 8'h19;
  picture_data[ 5199 ] = 8'h24;
  picture_data[ 5200 ] = 8'h00;
  picture_data[ 5201 ] = 8'hC2;
  picture_data[ 5202 ] = 8'h21;
  picture_data[ 5203 ] = 8'hC5;
  picture_data[ 5204 ] = 8'h21;
  picture_data[ 5205 ] = 8'hC5;
  picture_data[ 5206 ] = 8'h21;
  picture_data[ 5207 ] = 8'hC5;
  picture_data[ 5208 ] = 8'h19;
  picture_data[ 5209 ] = 8'h64;
  picture_data[ 5210 ] = 8'h19;
  picture_data[ 5211 ] = 8'h43;
  picture_data[ 5212 ] = 8'h08;
  picture_data[ 5213 ] = 8'hA1;
  picture_data[ 5214 ] = 8'h10;
  picture_data[ 5215 ] = 8'hA1;
  picture_data[ 5216 ] = 8'h21;
  picture_data[ 5217 ] = 8'h02;
  picture_data[ 5218 ] = 8'h10;
  picture_data[ 5219 ] = 8'hA1;
  picture_data[ 5220 ] = 8'h18;
  picture_data[ 5221 ] = 8'hE2;
  picture_data[ 5222 ] = 8'h18;
  picture_data[ 5223 ] = 8'hE1;
  picture_data[ 5224 ] = 8'h18;
  picture_data[ 5225 ] = 8'hE1;
  picture_data[ 5226 ] = 8'h19;
  picture_data[ 5227 ] = 8'h02;
  picture_data[ 5228 ] = 8'h19;
  picture_data[ 5229 ] = 8'h02;
  picture_data[ 5230 ] = 8'h18;
  picture_data[ 5231 ] = 8'hE1;
  picture_data[ 5232 ] = 8'h21;
  picture_data[ 5233 ] = 8'h42;
  picture_data[ 5234 ] = 8'h29;
  picture_data[ 5235 ] = 8'h83;
  picture_data[ 5236 ] = 8'h29;
  picture_data[ 5237 ] = 8'h43;
  picture_data[ 5238 ] = 8'h21;
  picture_data[ 5239 ] = 8'h23;
  picture_data[ 5240 ] = 8'h20;
  picture_data[ 5241 ] = 8'hC2;
  picture_data[ 5242 ] = 8'h29;
  picture_data[ 5243 ] = 8'h01;
  picture_data[ 5244 ] = 8'h39;
  picture_data[ 5245 ] = 8'h61;
  picture_data[ 5246 ] = 8'h41;
  picture_data[ 5247 ] = 8'h81;
  picture_data[ 5248 ] = 8'h39;
  picture_data[ 5249 ] = 8'h60;
  picture_data[ 5250 ] = 8'h41;
  picture_data[ 5251 ] = 8'hA0;
  picture_data[ 5252 ] = 8'h39;
  picture_data[ 5253 ] = 8'h61;
  picture_data[ 5254 ] = 8'h42;
  picture_data[ 5255 ] = 8'h04;
  picture_data[ 5256 ] = 8'h42;
  picture_data[ 5257 ] = 8'h25;
  picture_data[ 5258 ] = 8'h18;
  picture_data[ 5259 ] = 8'hE1;
  picture_data[ 5260 ] = 8'h19;
  picture_data[ 5261 ] = 8'h01;
  picture_data[ 5262 ] = 8'h19;
  picture_data[ 5263 ] = 8'h01;
  picture_data[ 5264 ] = 8'h19;
  picture_data[ 5265 ] = 8'h01;
  picture_data[ 5266 ] = 8'h18;
  picture_data[ 5267 ] = 8'hE1;
  picture_data[ 5268 ] = 8'h29;
  picture_data[ 5269 ] = 8'h63;
  picture_data[ 5270 ] = 8'h21;
  picture_data[ 5271 ] = 8'h42;
  picture_data[ 5272 ] = 8'h31;
  picture_data[ 5273 ] = 8'hA3;
  picture_data[ 5274 ] = 8'h3A;
  picture_data[ 5275 ] = 8'h05;
  picture_data[ 5276 ] = 8'h31;
  picture_data[ 5277 ] = 8'hA3;
  picture_data[ 5278 ] = 8'h31;
  picture_data[ 5279 ] = 8'hA3;
  picture_data[ 5280 ] = 8'h29;
  picture_data[ 5281 ] = 8'h83;
  picture_data[ 5282 ] = 8'h39;
  picture_data[ 5283 ] = 8'hC4;
  picture_data[ 5284 ] = 8'h21;
  picture_data[ 5285 ] = 8'h01;
  picture_data[ 5286 ] = 8'h31;
  picture_data[ 5287 ] = 8'hA3;
  picture_data[ 5288 ] = 8'h42;
  picture_data[ 5289 ] = 8'h05;
  picture_data[ 5290 ] = 8'h29;
  picture_data[ 5291 ] = 8'h63;
  picture_data[ 5292 ] = 8'h29;
  picture_data[ 5293 ] = 8'h62;
  picture_data[ 5294 ] = 8'h39;
  picture_data[ 5295 ] = 8'hC4;
  picture_data[ 5296 ] = 8'h31;
  picture_data[ 5297 ] = 8'h83;
  picture_data[ 5298 ] = 8'h29;
  picture_data[ 5299 ] = 8'h42;
  picture_data[ 5300 ] = 8'h42;
  picture_data[ 5301 ] = 8'h04;
  picture_data[ 5302 ] = 8'h4A;
  picture_data[ 5303 ] = 8'h24;
  picture_data[ 5304 ] = 8'h41;
  picture_data[ 5305 ] = 8'hC2;
  picture_data[ 5306 ] = 8'h39;
  picture_data[ 5307 ] = 8'hA2;
  picture_data[ 5308 ] = 8'h52;
  picture_data[ 5309 ] = 8'h44;
  picture_data[ 5310 ] = 8'h5A;
  picture_data[ 5311 ] = 8'h65;
  picture_data[ 5312 ] = 8'h49;
  picture_data[ 5313 ] = 8'hA2;
  picture_data[ 5314 ] = 8'h52;
  picture_data[ 5315 ] = 8'h04;
  picture_data[ 5316 ] = 8'h52;
  picture_data[ 5317 ] = 8'h05;
  picture_data[ 5318 ] = 8'h62;
  picture_data[ 5319 ] = 8'h66;
  picture_data[ 5320 ] = 8'h10;
  picture_data[ 5321 ] = 8'hA5;
  picture_data[ 5322 ] = 8'h00;
  picture_data[ 5323 ] = 8'h43;
  picture_data[ 5324 ] = 8'h08;
  picture_data[ 5325 ] = 8'hA4;
  picture_data[ 5326 ] = 8'h29;
  picture_data[ 5327 ] = 8'h88;
  picture_data[ 5328 ] = 8'h21;
  picture_data[ 5329 ] = 8'h47;
  picture_data[ 5330 ] = 8'h10;
  picture_data[ 5331 ] = 8'hE7;
  picture_data[ 5332 ] = 8'h10;
  picture_data[ 5333 ] = 8'hC7;
  picture_data[ 5334 ] = 8'h19;
  picture_data[ 5335 ] = 8'h07;
  picture_data[ 5336 ] = 8'h11;
  picture_data[ 5337 ] = 8'h05;
  picture_data[ 5338 ] = 8'h10;
  picture_data[ 5339 ] = 8'hE3;
  picture_data[ 5340 ] = 8'h08;
  picture_data[ 5341 ] = 8'hA2;
  picture_data[ 5342 ] = 8'h18;
  picture_data[ 5343 ] = 8'hE3;
  picture_data[ 5344 ] = 8'h08;
  picture_data[ 5345 ] = 8'h81;
  picture_data[ 5346 ] = 8'h18;
  picture_data[ 5347 ] = 8'hE3;
  picture_data[ 5348 ] = 8'h18;
  picture_data[ 5349 ] = 8'hE3;
  picture_data[ 5350 ] = 8'h08;
  picture_data[ 5351 ] = 8'hA2;
  picture_data[ 5352 ] = 8'h11;
  picture_data[ 5353 ] = 8'h23;
  picture_data[ 5354 ] = 8'h08;
  picture_data[ 5355 ] = 8'hC2;
  picture_data[ 5356 ] = 8'h19;
  picture_data[ 5357 ] = 8'h64;
  picture_data[ 5358 ] = 8'h21;
  picture_data[ 5359 ] = 8'h84;
  picture_data[ 5360 ] = 8'h11;
  picture_data[ 5361 ] = 8'h02;
  picture_data[ 5362 ] = 8'h21;
  picture_data[ 5363 ] = 8'h43;
  picture_data[ 5364 ] = 8'h10;
  picture_data[ 5365 ] = 8'hE1;
  picture_data[ 5366 ] = 8'h18;
  picture_data[ 5367 ] = 8'hE1;
  picture_data[ 5368 ] = 8'h18;
  picture_data[ 5369 ] = 8'hC1;
  picture_data[ 5370 ] = 8'h18;
  picture_data[ 5371 ] = 8'hC1;
  picture_data[ 5372 ] = 8'h18;
  picture_data[ 5373 ] = 8'hE1;
  picture_data[ 5374 ] = 8'h08;
  picture_data[ 5375 ] = 8'h80;
  picture_data[ 5376 ] = 8'h10;
  picture_data[ 5377 ] = 8'hC1;
  picture_data[ 5378 ] = 8'h21;
  picture_data[ 5379 ] = 8'h22;
  picture_data[ 5380 ] = 8'h18;
  picture_data[ 5381 ] = 8'hE2;
  picture_data[ 5382 ] = 8'h10;
  picture_data[ 5383 ] = 8'hE1;
  picture_data[ 5384 ] = 8'h19;
  picture_data[ 5385 ] = 8'h01;
  picture_data[ 5386 ] = 8'h19;
  picture_data[ 5387 ] = 8'h02;
  picture_data[ 5388 ] = 8'h29;
  picture_data[ 5389 ] = 8'hA5;
  picture_data[ 5390 ] = 8'h31;
  picture_data[ 5391 ] = 8'hA4;
  picture_data[ 5392 ] = 8'h18;
  picture_data[ 5393 ] = 8'hC0;
  picture_data[ 5394 ] = 8'h28;
  picture_data[ 5395 ] = 8'hE0;
  picture_data[ 5396 ] = 8'h51;
  picture_data[ 5397 ] = 8'hC1;
  picture_data[ 5398 ] = 8'h72;
  picture_data[ 5399 ] = 8'hC3;
  picture_data[ 5400 ] = 8'h83;
  picture_data[ 5401 ] = 8'h44;
  picture_data[ 5402 ] = 8'h62;
  picture_data[ 5403 ] = 8'h41;
  picture_data[ 5404 ] = 8'h39;
  picture_data[ 5405 ] = 8'h60;
  picture_data[ 5406 ] = 8'h41;
  picture_data[ 5407 ] = 8'hE2;
  picture_data[ 5408 ] = 8'h29;
  picture_data[ 5409 ] = 8'h62;
  picture_data[ 5410 ] = 8'h29;
  picture_data[ 5411 ] = 8'h62;
  picture_data[ 5412 ] = 8'h29;
  picture_data[ 5413 ] = 8'h63;
  picture_data[ 5414 ] = 8'h29;
  picture_data[ 5415 ] = 8'h63;
  picture_data[ 5416 ] = 8'h21;
  picture_data[ 5417 ] = 8'h42;
  picture_data[ 5418 ] = 8'h10;
  picture_data[ 5419 ] = 8'hA0;
  picture_data[ 5420 ] = 8'h21;
  picture_data[ 5421 ] = 8'h22;
  picture_data[ 5422 ] = 8'h29;
  picture_data[ 5423 ] = 8'h42;
  picture_data[ 5424 ] = 8'h31;
  picture_data[ 5425 ] = 8'h83;
  picture_data[ 5426 ] = 8'h31;
  picture_data[ 5427 ] = 8'h83;
  picture_data[ 5428 ] = 8'h29;
  picture_data[ 5429 ] = 8'h62;
  picture_data[ 5430 ] = 8'h29;
  picture_data[ 5431 ] = 8'h62;
  picture_data[ 5432 ] = 8'h31;
  picture_data[ 5433 ] = 8'h63;
  picture_data[ 5434 ] = 8'h31;
  picture_data[ 5435 ] = 8'hA3;
  picture_data[ 5436 ] = 8'h29;
  picture_data[ 5437 ] = 8'h62;
  picture_data[ 5438 ] = 8'h42;
  picture_data[ 5439 ] = 8'h05;
  picture_data[ 5440 ] = 8'h39;
  picture_data[ 5441 ] = 8'hC4;
  picture_data[ 5442 ] = 8'h10;
  picture_data[ 5443 ] = 8'hA0;
  picture_data[ 5444 ] = 8'h31;
  picture_data[ 5445 ] = 8'h63;
  picture_data[ 5446 ] = 8'h39;
  picture_data[ 5447 ] = 8'hE5;
  picture_data[ 5448 ] = 8'h29;
  picture_data[ 5449 ] = 8'h63;
  picture_data[ 5450 ] = 8'h39;
  picture_data[ 5451 ] = 8'hC4;
  picture_data[ 5452 ] = 8'h39;
  picture_data[ 5453 ] = 8'hE4;
  picture_data[ 5454 ] = 8'h42;
  picture_data[ 5455 ] = 8'h24;
  picture_data[ 5456 ] = 8'h4A;
  picture_data[ 5457 ] = 8'h24;
  picture_data[ 5458 ] = 8'h41;
  picture_data[ 5459 ] = 8'hE3;
  picture_data[ 5460 ] = 8'h39;
  picture_data[ 5461 ] = 8'h81;
  picture_data[ 5462 ] = 8'h52;
  picture_data[ 5463 ] = 8'h65;
  picture_data[ 5464 ] = 8'h39;
  picture_data[ 5465 ] = 8'h62;
  picture_data[ 5466 ] = 8'h52;
  picture_data[ 5467 ] = 8'h25;
  picture_data[ 5468 ] = 8'h52;
  picture_data[ 5469 ] = 8'h26;
  picture_data[ 5470 ] = 8'h52;
  picture_data[ 5471 ] = 8'h46;
  picture_data[ 5472 ] = 8'h00;
  picture_data[ 5473 ] = 8'h65;
  picture_data[ 5474 ] = 8'h00;
  picture_data[ 5475 ] = 8'h85;
  picture_data[ 5476 ] = 8'h08;
  picture_data[ 5477 ] = 8'hA6;
  picture_data[ 5478 ] = 8'h21;
  picture_data[ 5479 ] = 8'h8B;
  picture_data[ 5480 ] = 8'h11;
  picture_data[ 5481 ] = 8'h2A;
  picture_data[ 5482 ] = 8'h08;
  picture_data[ 5483 ] = 8'hE9;
  picture_data[ 5484 ] = 8'h08;
  picture_data[ 5485 ] = 8'hCA;
  picture_data[ 5486 ] = 8'h29;
  picture_data[ 5487 ] = 8'hAC;
  picture_data[ 5488 ] = 8'h19;
  picture_data[ 5489 ] = 8'h48;
  picture_data[ 5490 ] = 8'h00;
  picture_data[ 5491 ] = 8'h82;
  picture_data[ 5492 ] = 8'h10;
  picture_data[ 5493 ] = 8'hE3;
  picture_data[ 5494 ] = 8'h10;
  picture_data[ 5495 ] = 8'hE2;
  picture_data[ 5496 ] = 8'h10;
  picture_data[ 5497 ] = 8'hC2;
  picture_data[ 5498 ] = 8'h10;
  picture_data[ 5499 ] = 8'hC1;
  picture_data[ 5500 ] = 8'h10;
  picture_data[ 5501 ] = 8'hA1;
  picture_data[ 5502 ] = 8'h18;
  picture_data[ 5503 ] = 8'hE2;
  picture_data[ 5504 ] = 8'h08;
  picture_data[ 5505 ] = 8'hC2;
  picture_data[ 5506 ] = 8'h21;
  picture_data[ 5507 ] = 8'h64;
  picture_data[ 5508 ] = 8'h31;
  picture_data[ 5509 ] = 8'hC6;
  picture_data[ 5510 ] = 8'h10;
  picture_data[ 5511 ] = 8'hE2;
  picture_data[ 5512 ] = 8'h10;
  picture_data[ 5513 ] = 8'hC1;
  picture_data[ 5514 ] = 8'h10;
  picture_data[ 5515 ] = 8'hA1;
  picture_data[ 5516 ] = 8'h19;
  picture_data[ 5517 ] = 8'h02;
  picture_data[ 5518 ] = 8'h10;
  picture_data[ 5519 ] = 8'hA1;
  picture_data[ 5520 ] = 8'h18;
  picture_data[ 5521 ] = 8'hC1;
  picture_data[ 5522 ] = 8'h10;
  picture_data[ 5523 ] = 8'hA0;
  picture_data[ 5524 ] = 8'h19;
  picture_data[ 5525 ] = 8'h02;
  picture_data[ 5526 ] = 8'h18;
  picture_data[ 5527 ] = 8'hE1;
  picture_data[ 5528 ] = 8'h08;
  picture_data[ 5529 ] = 8'h60;
  picture_data[ 5530 ] = 8'h10;
  picture_data[ 5531 ] = 8'hC1;
  picture_data[ 5532 ] = 8'h10;
  picture_data[ 5533 ] = 8'hE1;
  picture_data[ 5534 ] = 8'h10;
  picture_data[ 5535 ] = 8'hC1;
  picture_data[ 5536 ] = 8'h10;
  picture_data[ 5537 ] = 8'hC1;
  picture_data[ 5538 ] = 8'h19;
  picture_data[ 5539 ] = 8'h02;
  picture_data[ 5540 ] = 8'h19;
  picture_data[ 5541 ] = 8'h43;
  picture_data[ 5542 ] = 8'h19;
  picture_data[ 5543 ] = 8'h22;
  picture_data[ 5544 ] = 8'h21;
  picture_data[ 5545 ] = 8'h20;
  picture_data[ 5546 ] = 8'h41;
  picture_data[ 5547 ] = 8'hA0;
  picture_data[ 5548 ] = 8'h6A;
  picture_data[ 5549 ] = 8'hA2;
  picture_data[ 5550 ] = 8'hD5;
  picture_data[ 5551 ] = 8'hCC;
  picture_data[ 5552 ] = 8'hFF;
  picture_data[ 5553 ] = 8'h52;
  picture_data[ 5554 ] = 8'hC5;
  picture_data[ 5555 ] = 8'h2A;
  picture_data[ 5556 ] = 8'h6A;
  picture_data[ 5557 ] = 8'hE3;
  picture_data[ 5558 ] = 8'h52;
  picture_data[ 5559 ] = 8'h63;
  picture_data[ 5560 ] = 8'h31;
  picture_data[ 5561 ] = 8'h82;
  picture_data[ 5562 ] = 8'h21;
  picture_data[ 5563 ] = 8'h21;
  picture_data[ 5564 ] = 8'h21;
  picture_data[ 5565 ] = 8'h22;
  picture_data[ 5566 ] = 8'h29;
  picture_data[ 5567 ] = 8'h42;
  picture_data[ 5568 ] = 8'h21;
  picture_data[ 5569 ] = 8'h02;
  picture_data[ 5570 ] = 8'h21;
  picture_data[ 5571 ] = 8'h22;
  picture_data[ 5572 ] = 8'h29;
  picture_data[ 5573 ] = 8'h42;
  picture_data[ 5574 ] = 8'h29;
  picture_data[ 5575 ] = 8'h22;
  picture_data[ 5576 ] = 8'h31;
  picture_data[ 5577 ] = 8'hA3;
  picture_data[ 5578 ] = 8'h31;
  picture_data[ 5579 ] = 8'h63;
  picture_data[ 5580 ] = 8'h29;
  picture_data[ 5581 ] = 8'h21;
  picture_data[ 5582 ] = 8'h29;
  picture_data[ 5583 ] = 8'h21;
  picture_data[ 5584 ] = 8'h31;
  picture_data[ 5585 ] = 8'h83;
  picture_data[ 5586 ] = 8'h31;
  picture_data[ 5587 ] = 8'h82;
  picture_data[ 5588 ] = 8'h31;
  picture_data[ 5589 ] = 8'h83;
  picture_data[ 5590 ] = 8'h39;
  picture_data[ 5591 ] = 8'hC4;
  picture_data[ 5592 ] = 8'h39;
  picture_data[ 5593 ] = 8'hE5;
  picture_data[ 5594 ] = 8'h21;
  picture_data[ 5595 ] = 8'h01;
  picture_data[ 5596 ] = 8'h31;
  picture_data[ 5597 ] = 8'hA4;
  picture_data[ 5598 ] = 8'h31;
  picture_data[ 5599 ] = 8'hA4;
  picture_data[ 5600 ] = 8'h31;
  picture_data[ 5601 ] = 8'hA3;
  picture_data[ 5602 ] = 8'h39;
  picture_data[ 5603 ] = 8'hE4;
  picture_data[ 5604 ] = 8'h39;
  picture_data[ 5605 ] = 8'hC3;
  picture_data[ 5606 ] = 8'h31;
  picture_data[ 5607 ] = 8'hA3;
  picture_data[ 5608 ] = 8'h39;
  picture_data[ 5609 ] = 8'hA3;
  picture_data[ 5610 ] = 8'h31;
  picture_data[ 5611 ] = 8'h82;
  picture_data[ 5612 ] = 8'h31;
  picture_data[ 5613 ] = 8'h62;
  picture_data[ 5614 ] = 8'h52;
  picture_data[ 5615 ] = 8'h66;
  picture_data[ 5616 ] = 8'h41;
  picture_data[ 5617 ] = 8'hC4;
  picture_data[ 5618 ] = 8'h4A;
  picture_data[ 5619 ] = 8'h26;
  picture_data[ 5620 ] = 8'h41;
  picture_data[ 5621 ] = 8'hE5;
  picture_data[ 5622 ] = 8'h41;
  picture_data[ 5623 ] = 8'hE5;
  picture_data[ 5624 ] = 8'h66;
  picture_data[ 5625 ] = 8'h00;
  picture_data[ 5626 ] = 8'h88;
  picture_data[ 5627 ] = 8'h09;
  picture_data[ 5628 ] = 8'h0B;
  picture_data[ 5629 ] = 8'h19;
  picture_data[ 5630 ] = 8'hD0;
  picture_data[ 5631 ] = 8'h09;
  picture_data[ 5632 ] = 8'h4F;
  picture_data[ 5633 ] = 8'h09;
  picture_data[ 5634 ] = 8'h0F;
  picture_data[ 5635 ] = 8'h00;
  picture_data[ 5636 ] = 8'hCE;
  picture_data[ 5637 ] = 8'h11;
  picture_data[ 5638 ] = 8'h0C;
  picture_data[ 5639 ] = 8'h21;
  picture_data[ 5640 ] = 8'h8A;
  picture_data[ 5641 ] = 8'h19;
  picture_data[ 5642 ] = 8'h26;
  picture_data[ 5643 ] = 8'h10;
  picture_data[ 5644 ] = 8'hC3;
  picture_data[ 5645 ] = 8'h10;
  picture_data[ 5646 ] = 8'hE3;
  picture_data[ 5647 ] = 8'h10;
  picture_data[ 5648 ] = 8'hE2;
  picture_data[ 5649 ] = 8'h10;
  picture_data[ 5650 ] = 8'hC2;
  picture_data[ 5651 ] = 8'h08;
  picture_data[ 5652 ] = 8'hA1;
  picture_data[ 5653 ] = 8'h18;
  picture_data[ 5654 ] = 8'hE2;
  picture_data[ 5655 ] = 8'h10;
  picture_data[ 5656 ] = 8'hA1;
  picture_data[ 5657 ] = 8'h19;
  picture_data[ 5658 ] = 8'h03;
  picture_data[ 5659 ] = 8'h18;
  picture_data[ 5660 ] = 8'hE2;
  picture_data[ 5661 ] = 8'h19;
  picture_data[ 5662 ] = 8'h03;
  picture_data[ 5663 ] = 8'h21;
  picture_data[ 5664 ] = 8'h23;
  picture_data[ 5665 ] = 8'h18;
  picture_data[ 5666 ] = 8'hE2;
  picture_data[ 5667 ] = 8'h10;
  picture_data[ 5668 ] = 8'hC1;
  picture_data[ 5669 ] = 8'h19;
  picture_data[ 5670 ] = 8'h02;
  picture_data[ 5671 ] = 8'h19;
  picture_data[ 5672 ] = 8'h02;
  picture_data[ 5673 ] = 8'h18;
  picture_data[ 5674 ] = 8'hE1;
  picture_data[ 5675 ] = 8'h18;
  picture_data[ 5676 ] = 8'hE1;
  picture_data[ 5677 ] = 8'h21;
  picture_data[ 5678 ] = 8'h22;
  picture_data[ 5679 ] = 8'h18;
  picture_data[ 5680 ] = 8'hE1;
  picture_data[ 5681 ] = 8'h10;
  picture_data[ 5682 ] = 8'hA1;
  picture_data[ 5683 ] = 8'h10;
  picture_data[ 5684 ] = 8'hA0;
  picture_data[ 5685 ] = 8'h08;
  picture_data[ 5686 ] = 8'hA0;
  picture_data[ 5687 ] = 8'h10;
  picture_data[ 5688 ] = 8'hA1;
  picture_data[ 5689 ] = 8'h19;
  picture_data[ 5690 ] = 8'h02;
  picture_data[ 5691 ] = 8'h10;
  picture_data[ 5692 ] = 8'hE2;
  picture_data[ 5693 ] = 8'h19;
  picture_data[ 5694 ] = 8'h02;
  picture_data[ 5695 ] = 8'h29;
  picture_data[ 5696 ] = 8'h62;
  picture_data[ 5697 ] = 8'h39;
  picture_data[ 5698 ] = 8'h80;
  picture_data[ 5699 ] = 8'h49;
  picture_data[ 5700 ] = 8'h80;
  picture_data[ 5701 ] = 8'h9C;
  picture_data[ 5702 ] = 8'h05;
  picture_data[ 5703 ] = 8'hF6;
  picture_data[ 5704 ] = 8'hAF;
  picture_data[ 5705 ] = 8'hCD;
  picture_data[ 5706 ] = 8'hAC;
  picture_data[ 5707 ] = 8'h83;
  picture_data[ 5708 ] = 8'h86;
  picture_data[ 5709 ] = 8'h52;
  picture_data[ 5710 ] = 8'h43;
  picture_data[ 5711 ] = 8'h42;
  picture_data[ 5712 ] = 8'h04;
  picture_data[ 5713 ] = 8'h29;
  picture_data[ 5714 ] = 8'h42;
  picture_data[ 5715 ] = 8'h31;
  picture_data[ 5716 ] = 8'h63;
  picture_data[ 5717 ] = 8'h21;
  picture_data[ 5718 ] = 8'h01;
  picture_data[ 5719 ] = 8'h20;
  picture_data[ 5720 ] = 8'hE1;
  picture_data[ 5721 ] = 8'h21;
  picture_data[ 5722 ] = 8'h02;
  picture_data[ 5723 ] = 8'h29;
  picture_data[ 5724 ] = 8'h22;
  picture_data[ 5725 ] = 8'h29;
  picture_data[ 5726 ] = 8'h42;
  picture_data[ 5727 ] = 8'h31;
  picture_data[ 5728 ] = 8'h63;
  picture_data[ 5729 ] = 8'h31;
  picture_data[ 5730 ] = 8'h62;
  picture_data[ 5731 ] = 8'h31;
  picture_data[ 5732 ] = 8'h62;
  picture_data[ 5733 ] = 8'h29;
  picture_data[ 5734 ] = 8'h21;
  picture_data[ 5735 ] = 8'h29;
  picture_data[ 5736 ] = 8'h41;
  picture_data[ 5737 ] = 8'h31;
  picture_data[ 5738 ] = 8'h62;
  picture_data[ 5739 ] = 8'h29;
  picture_data[ 5740 ] = 8'h41;
  picture_data[ 5741 ] = 8'h29;
  picture_data[ 5742 ] = 8'h22;
  picture_data[ 5743 ] = 8'h39;
  picture_data[ 5744 ] = 8'hC4;
  picture_data[ 5745 ] = 8'h39;
  picture_data[ 5746 ] = 8'hC4;
  picture_data[ 5747 ] = 8'h29;
  picture_data[ 5748 ] = 8'h63;
  picture_data[ 5749 ] = 8'h29;
  picture_data[ 5750 ] = 8'h63;
  picture_data[ 5751 ] = 8'h39;
  picture_data[ 5752 ] = 8'hE5;
  picture_data[ 5753 ] = 8'h39;
  picture_data[ 5754 ] = 8'hC4;
  picture_data[ 5755 ] = 8'h42;
  picture_data[ 5756 ] = 8'h05;
  picture_data[ 5757 ] = 8'h39;
  picture_data[ 5758 ] = 8'hC4;
  picture_data[ 5759 ] = 8'h31;
  picture_data[ 5760 ] = 8'hA3;
  picture_data[ 5761 ] = 8'h39;
  picture_data[ 5762 ] = 8'hC4;
  picture_data[ 5763 ] = 8'h42;
  picture_data[ 5764 ] = 8'h05;
  picture_data[ 5765 ] = 8'h39;
  picture_data[ 5766 ] = 8'hA4;
  picture_data[ 5767 ] = 8'h4A;
  picture_data[ 5768 ] = 8'h26;
  picture_data[ 5769 ] = 8'h41;
  picture_data[ 5770 ] = 8'hE5;
  picture_data[ 5771 ] = 8'h29;
  picture_data[ 5772 ] = 8'h43;
  picture_data[ 5773 ] = 8'h29;
  picture_data[ 5774 ] = 8'h43;
  picture_data[ 5775 ] = 8'h49;
  picture_data[ 5776 ] = 8'h00;
  picture_data[ 5777 ] = 8'hAC;
  picture_data[ 5778 ] = 8'h00;
  picture_data[ 5779 ] = 8'hF0;
  picture_data[ 5780 ] = 8'h01;
  picture_data[ 5781 ] = 8'h75;
  picture_data[ 5782 ] = 8'h09;
  picture_data[ 5783 ] = 8'hD8;
  picture_data[ 5784 ] = 8'h01;
  picture_data[ 5785 ] = 8'h97;
  picture_data[ 5786 ] = 8'h00;
  picture_data[ 5787 ] = 8'hF3;
  picture_data[ 5788 ] = 8'h11;
  picture_data[ 5789 ] = 8'h30;
  picture_data[ 5790 ] = 8'h10;
  picture_data[ 5791 ] = 8'hEA;
  picture_data[ 5792 ] = 8'h29;
  picture_data[ 5793 ] = 8'h89;
  picture_data[ 5794 ] = 8'h10;
  picture_data[ 5795 ] = 8'hE5;
  picture_data[ 5796 ] = 8'h19;
  picture_data[ 5797 ] = 8'h05;
  picture_data[ 5798 ] = 8'h00;
  picture_data[ 5799 ] = 8'h82;
  picture_data[ 5800 ] = 8'h00;
  picture_data[ 5801 ] = 8'h81;
  picture_data[ 5802 ] = 8'h10;
  picture_data[ 5803 ] = 8'hA1;
  picture_data[ 5804 ] = 8'h18;
  picture_data[ 5805 ] = 8'hC1;
  picture_data[ 5806 ] = 8'h10;
  picture_data[ 5807 ] = 8'h81;
  picture_data[ 5808 ] = 8'h18;
  picture_data[ 5809 ] = 8'hC2;
  picture_data[ 5810 ] = 8'h21;
  picture_data[ 5811 ] = 8'h03;
  picture_data[ 5812 ] = 8'h10;
  picture_data[ 5813 ] = 8'h81;
  picture_data[ 5814 ] = 8'h08;
  picture_data[ 5815 ] = 8'h80;
  picture_data[ 5816 ] = 8'h10;
  picture_data[ 5817 ] = 8'hA0;
  picture_data[ 5818 ] = 8'h10;
  picture_data[ 5819 ] = 8'hC1;
  picture_data[ 5820 ] = 8'h10;
  picture_data[ 5821 ] = 8'hC1;
  picture_data[ 5822 ] = 8'h18;
  picture_data[ 5823 ] = 8'hE2;
  picture_data[ 5824 ] = 8'h29;
  picture_data[ 5825 ] = 8'h63;
  picture_data[ 5826 ] = 8'h08;
  picture_data[ 5827 ] = 8'h80;
  picture_data[ 5828 ] = 8'h10;
  picture_data[ 5829 ] = 8'hA1;
  picture_data[ 5830 ] = 8'h21;
  picture_data[ 5831 ] = 8'h43;
  picture_data[ 5832 ] = 8'h18;
  picture_data[ 5833 ] = 8'hE1;
  picture_data[ 5834 ] = 8'h00;
  picture_data[ 5835 ] = 8'h40;
  picture_data[ 5836 ] = 8'h10;
  picture_data[ 5837 ] = 8'hC1;
  picture_data[ 5838 ] = 8'h10;
  picture_data[ 5839 ] = 8'h80;
  picture_data[ 5840 ] = 8'h10;
  picture_data[ 5841 ] = 8'h81;
  picture_data[ 5842 ] = 8'h19;
  picture_data[ 5843 ] = 8'h03;
  picture_data[ 5844 ] = 8'h10;
  picture_data[ 5845 ] = 8'hA1;
  picture_data[ 5846 ] = 8'h29;
  picture_data[ 5847 ] = 8'h22;
  picture_data[ 5848 ] = 8'h18;
  picture_data[ 5849 ] = 8'hA0;
  picture_data[ 5850 ] = 8'h41;
  picture_data[ 5851 ] = 8'h80;
  picture_data[ 5852 ] = 8'h5A;
  picture_data[ 5853 ] = 8'h00;
  picture_data[ 5854 ] = 8'h83;
  picture_data[ 5855 ] = 8'h45;
  picture_data[ 5856 ] = 8'h73;
  picture_data[ 5857 ] = 8'h04;
  picture_data[ 5858 ] = 8'h41;
  picture_data[ 5859 ] = 8'hA0;
  picture_data[ 5860 ] = 8'h39;
  picture_data[ 5861 ] = 8'hA2;
  picture_data[ 5862 ] = 8'h39;
  picture_data[ 5863 ] = 8'hA3;
  picture_data[ 5864 ] = 8'h31;
  picture_data[ 5865 ] = 8'h63;
  picture_data[ 5866 ] = 8'h29;
  picture_data[ 5867 ] = 8'h22;
  picture_data[ 5868 ] = 8'h31;
  picture_data[ 5869 ] = 8'h43;
  picture_data[ 5870 ] = 8'h29;
  picture_data[ 5871 ] = 8'h23;
  picture_data[ 5872 ] = 8'h18;
  picture_data[ 5873 ] = 8'hC1;
  picture_data[ 5874 ] = 8'h29;
  picture_data[ 5875 ] = 8'h22;
  picture_data[ 5876 ] = 8'h31;
  picture_data[ 5877 ] = 8'h83;
  picture_data[ 5878 ] = 8'h29;
  picture_data[ 5879 ] = 8'h42;
  picture_data[ 5880 ] = 8'h31;
  picture_data[ 5881 ] = 8'h83;
  picture_data[ 5882 ] = 8'h31;
  picture_data[ 5883 ] = 8'h83;
  picture_data[ 5884 ] = 8'h29;
  picture_data[ 5885 ] = 8'h41;
  picture_data[ 5886 ] = 8'h31;
  picture_data[ 5887 ] = 8'h42;
  picture_data[ 5888 ] = 8'h29;
  picture_data[ 5889 ] = 8'h42;
  picture_data[ 5890 ] = 8'h39;
  picture_data[ 5891 ] = 8'hA3;
  picture_data[ 5892 ] = 8'h31;
  picture_data[ 5893 ] = 8'hA3;
  picture_data[ 5894 ] = 8'h29;
  picture_data[ 5895 ] = 8'h42;
  picture_data[ 5896 ] = 8'h31;
  picture_data[ 5897 ] = 8'h83;
  picture_data[ 5898 ] = 8'h31;
  picture_data[ 5899 ] = 8'h83;
  picture_data[ 5900 ] = 8'h29;
  picture_data[ 5901 ] = 8'h63;
  picture_data[ 5902 ] = 8'h31;
  picture_data[ 5903 ] = 8'h83;
  picture_data[ 5904 ] = 8'h31;
  picture_data[ 5905 ] = 8'h82;
  picture_data[ 5906 ] = 8'h31;
  picture_data[ 5907 ] = 8'h83;
  picture_data[ 5908 ] = 8'h39;
  picture_data[ 5909 ] = 8'hC4;
  picture_data[ 5910 ] = 8'h41;
  picture_data[ 5911 ] = 8'hE5;
  picture_data[ 5912 ] = 8'h31;
  picture_data[ 5913 ] = 8'h83;
  picture_data[ 5914 ] = 8'h4A;
  picture_data[ 5915 ] = 8'h26;
  picture_data[ 5916 ] = 8'h63;
  picture_data[ 5917 ] = 8'h0A;
  picture_data[ 5918 ] = 8'h31;
  picture_data[ 5919 ] = 8'h84;
  picture_data[ 5920 ] = 8'h31;
  picture_data[ 5921 ] = 8'h84;
  picture_data[ 5922 ] = 8'h20;
  picture_data[ 5923 ] = 8'hE2;
  picture_data[ 5924 ] = 8'h18;
  picture_data[ 5925 ] = 8'hC1;
  picture_data[ 5926 ] = 8'h08;
  picture_data[ 5927 ] = 8'h8A;
  picture_data[ 5928 ] = 8'h00;
  picture_data[ 5929 ] = 8'h6C;
  picture_data[ 5930 ] = 8'h09;
  picture_data[ 5931 ] = 8'h75;
  picture_data[ 5932 ] = 8'h1A;
  picture_data[ 5933 ] = 8'h7B;
  picture_data[ 5934 ] = 8'h22;
  picture_data[ 5935 ] = 8'hDF;
  picture_data[ 5936 ] = 8'h12;
  picture_data[ 5937 ] = 8'h3C;
  picture_data[ 5938 ] = 8'h11;
  picture_data[ 5939 ] = 8'h97;
  picture_data[ 5940 ] = 8'h00;
  picture_data[ 5941 ] = 8'hD0;
  picture_data[ 5942 ] = 8'h19;
  picture_data[ 5943 ] = 8'h4C;
  picture_data[ 5944 ] = 8'h19;
  picture_data[ 5945 ] = 8'h08;
  picture_data[ 5946 ] = 8'h21;
  picture_data[ 5947 ] = 8'h48;
  picture_data[ 5948 ] = 8'h19;
  picture_data[ 5949 ] = 8'h26;
  picture_data[ 5950 ] = 8'h08;
  picture_data[ 5951 ] = 8'hA4;
  picture_data[ 5952 ] = 8'h08;
  picture_data[ 5953 ] = 8'hA2;
  picture_data[ 5954 ] = 8'h08;
  picture_data[ 5955 ] = 8'h81;
  picture_data[ 5956 ] = 8'h08;
  picture_data[ 5957 ] = 8'h60;
  picture_data[ 5958 ] = 8'h08;
  picture_data[ 5959 ] = 8'h61;
  picture_data[ 5960 ] = 8'h10;
  picture_data[ 5961 ] = 8'hA1;
  picture_data[ 5962 ] = 8'h08;
  picture_data[ 5963 ] = 8'h61;
  picture_data[ 5964 ] = 8'h10;
  picture_data[ 5965 ] = 8'h81;
  picture_data[ 5966 ] = 8'h18;
  picture_data[ 5967 ] = 8'hC2;
  picture_data[ 5968 ] = 8'h18;
  picture_data[ 5969 ] = 8'hE2;
  picture_data[ 5970 ] = 8'h18;
  picture_data[ 5971 ] = 8'hC2;
  picture_data[ 5972 ] = 8'h08;
  picture_data[ 5973 ] = 8'h60;
  picture_data[ 5974 ] = 8'h19;
  picture_data[ 5975 ] = 8'h02;
  picture_data[ 5976 ] = 8'h18;
  picture_data[ 5977 ] = 8'hC2;
  picture_data[ 5978 ] = 8'h08;
  picture_data[ 5979 ] = 8'h60;
  picture_data[ 5980 ] = 8'h10;
  picture_data[ 5981 ] = 8'hC1;
  picture_data[ 5982 ] = 8'h08;
  picture_data[ 5983 ] = 8'h60;
  picture_data[ 5984 ] = 8'h10;
  picture_data[ 5985 ] = 8'hA1;
  picture_data[ 5986 ] = 8'h21;
  picture_data[ 5987 ] = 8'h02;
  picture_data[ 5988 ] = 8'h10;
  picture_data[ 5989 ] = 8'h80;
  picture_data[ 5990 ] = 8'h10;
  picture_data[ 5991 ] = 8'h81;
  picture_data[ 5992 ] = 8'h18;
  picture_data[ 5993 ] = 8'hC2;
  picture_data[ 5994 ] = 8'h18;
  picture_data[ 5995 ] = 8'hC2;
  picture_data[ 5996 ] = 8'h18;
  picture_data[ 5997 ] = 8'hC2;
  picture_data[ 5998 ] = 8'h10;
  picture_data[ 5999 ] = 8'h80;
  picture_data[ 6000 ] = 8'h10;
  picture_data[ 6001 ] = 8'h80;
  picture_data[ 6002 ] = 8'h39;
  picture_data[ 6003 ] = 8'h82;
  picture_data[ 6004 ] = 8'h28;
  picture_data[ 6005 ] = 8'hE0;
  picture_data[ 6006 ] = 8'h31;
  picture_data[ 6007 ] = 8'h00;
  picture_data[ 6008 ] = 8'h39;
  picture_data[ 6009 ] = 8'h40;
  picture_data[ 6010 ] = 8'h41;
  picture_data[ 6011 ] = 8'hC3;
  picture_data[ 6012 ] = 8'h29;
  picture_data[ 6013 ] = 8'h21;
  picture_data[ 6014 ] = 8'h29;
  picture_data[ 6015 ] = 8'h22;
  picture_data[ 6016 ] = 8'h29;
  picture_data[ 6017 ] = 8'h02;
  picture_data[ 6018 ] = 8'h31;
  picture_data[ 6019 ] = 8'h23;
  picture_data[ 6020 ] = 8'h31;
  picture_data[ 6021 ] = 8'h43;
  picture_data[ 6022 ] = 8'h29;
  picture_data[ 6023 ] = 8'h23;
  picture_data[ 6024 ] = 8'h20;
  picture_data[ 6025 ] = 8'hE2;
  picture_data[ 6026 ] = 8'h21;
  picture_data[ 6027 ] = 8'h22;
  picture_data[ 6028 ] = 8'h21;
  picture_data[ 6029 ] = 8'h22;
  picture_data[ 6030 ] = 8'h29;
  picture_data[ 6031 ] = 8'h22;
  picture_data[ 6032 ] = 8'h39;
  picture_data[ 6033 ] = 8'hA4;
  picture_data[ 6034 ] = 8'h29;
  picture_data[ 6035 ] = 8'h42;
  picture_data[ 6036 ] = 8'h31;
  picture_data[ 6037 ] = 8'h62;
  picture_data[ 6038 ] = 8'h39;
  picture_data[ 6039 ] = 8'hA2;
  picture_data[ 6040 ] = 8'h31;
  picture_data[ 6041 ] = 8'h62;
  picture_data[ 6042 ] = 8'h29;
  picture_data[ 6043 ] = 8'h41;
  picture_data[ 6044 ] = 8'h31;
  picture_data[ 6045 ] = 8'h62;
  picture_data[ 6046 ] = 8'h31;
  picture_data[ 6047 ] = 8'hA3;
  picture_data[ 6048 ] = 8'h31;
  picture_data[ 6049 ] = 8'hA3;
  picture_data[ 6050 ] = 8'h31;
  picture_data[ 6051 ] = 8'h83;
  picture_data[ 6052 ] = 8'h39;
  picture_data[ 6053 ] = 8'hA4;
  picture_data[ 6054 ] = 8'h29;
  picture_data[ 6055 ] = 8'h62;
  picture_data[ 6056 ] = 8'h42;
  picture_data[ 6057 ] = 8'h04;
  picture_data[ 6058 ] = 8'h41;
  picture_data[ 6059 ] = 8'hE5;
  picture_data[ 6060 ] = 8'h42;
  picture_data[ 6061 ] = 8'h25;
  picture_data[ 6062 ] = 8'h41;
  picture_data[ 6063 ] = 8'hE5;
  picture_data[ 6064 ] = 8'h41;
  picture_data[ 6065 ] = 8'hE5;
  picture_data[ 6066 ] = 8'h39;
  picture_data[ 6067 ] = 8'hC5;
  picture_data[ 6068 ] = 8'h39;
  picture_data[ 6069 ] = 8'hA5;
  picture_data[ 6070 ] = 8'h10;
  picture_data[ 6071 ] = 8'h81;
  picture_data[ 6072 ] = 8'h31;
  picture_data[ 6073 ] = 8'h64;
  picture_data[ 6074 ] = 8'h31;
  picture_data[ 6075 ] = 8'h64;
  picture_data[ 6076 ] = 8'h21;
  picture_data[ 6077 ] = 8'h02;
  picture_data[ 6078 ] = 8'h08;
  picture_data[ 6079 ] = 8'hC9;
  picture_data[ 6080 ] = 8'h00;
  picture_data[ 6081 ] = 8'h8B;
  picture_data[ 6082 ] = 8'h11;
  picture_data[ 6083 ] = 8'hF5;
  picture_data[ 6084 ] = 8'h12;
  picture_data[ 6085 ] = 8'h5A;
  picture_data[ 6086 ] = 8'h12;
  picture_data[ 6087 ] = 8'h5C;
  picture_data[ 6088 ] = 8'h2A;
  picture_data[ 6089 ] = 8'hFE;
  picture_data[ 6090 ] = 8'h09;
  picture_data[ 6091 ] = 8'h96;
  picture_data[ 6092 ] = 8'h00;
  picture_data[ 6093 ] = 8'hCF;
  picture_data[ 6094 ] = 8'h19;
  picture_data[ 6095 ] = 8'h2B;
  picture_data[ 6096 ] = 8'h19;
  picture_data[ 6097 ] = 8'h07;
  picture_data[ 6098 ] = 8'h19;
  picture_data[ 6099 ] = 8'h28;
  picture_data[ 6100 ] = 8'h10;
  picture_data[ 6101 ] = 8'hA6;
  picture_data[ 6102 ] = 8'h10;
  picture_data[ 6103 ] = 8'hE7;
  picture_data[ 6104 ] = 8'h08;
  picture_data[ 6105 ] = 8'hA5;
  picture_data[ 6106 ] = 8'h08;
  picture_data[ 6107 ] = 8'h83;
  picture_data[ 6108 ] = 8'h10;
  picture_data[ 6109 ] = 8'h82;
  picture_data[ 6110 ] = 8'h08;
  picture_data[ 6111 ] = 8'h81;
  picture_data[ 6112 ] = 8'h10;
  picture_data[ 6113 ] = 8'hA2;
  picture_data[ 6114 ] = 8'h08;
  picture_data[ 6115 ] = 8'h81;
  picture_data[ 6116 ] = 8'h08;
  picture_data[ 6117 ] = 8'h81;
  picture_data[ 6118 ] = 8'h10;
  picture_data[ 6119 ] = 8'hC2;
  picture_data[ 6120 ] = 8'h10;
  picture_data[ 6121 ] = 8'hA1;
  picture_data[ 6122 ] = 8'h08;
  picture_data[ 6123 ] = 8'h81;
  picture_data[ 6124 ] = 8'h10;
  picture_data[ 6125 ] = 8'hC1;
  picture_data[ 6126 ] = 8'h10;
  picture_data[ 6127 ] = 8'hA1;
  picture_data[ 6128 ] = 8'h10;
  picture_data[ 6129 ] = 8'hA1;
  picture_data[ 6130 ] = 8'h08;
  picture_data[ 6131 ] = 8'h81;
  picture_data[ 6132 ] = 8'h08;
  picture_data[ 6133 ] = 8'h81;
  picture_data[ 6134 ] = 8'h10;
  picture_data[ 6135 ] = 8'h81;
  picture_data[ 6136 ] = 8'h10;
  picture_data[ 6137 ] = 8'h81;
  picture_data[ 6138 ] = 8'h10;
  picture_data[ 6139 ] = 8'hA1;
  picture_data[ 6140 ] = 8'h18;
  picture_data[ 6141 ] = 8'hE2;
  picture_data[ 6142 ] = 8'h18;
  picture_data[ 6143 ] = 8'hA1;
  picture_data[ 6144 ] = 8'h10;
  picture_data[ 6145 ] = 8'h81;
  picture_data[ 6146 ] = 8'h20;
  picture_data[ 6147 ] = 8'hE2;
  picture_data[ 6148 ] = 8'h18;
  picture_data[ 6149 ] = 8'hC2;
  picture_data[ 6150 ] = 8'h10;
  picture_data[ 6151 ] = 8'h81;
  picture_data[ 6152 ] = 8'h18;
  picture_data[ 6153 ] = 8'hE1;
  picture_data[ 6154 ] = 8'h21;
  picture_data[ 6155 ] = 8'h02;
  picture_data[ 6156 ] = 8'h29;
  picture_data[ 6157 ] = 8'h02;
  picture_data[ 6158 ] = 8'h20;
  picture_data[ 6159 ] = 8'hC0;
  picture_data[ 6160 ] = 8'h29;
  picture_data[ 6161 ] = 8'h01;
  picture_data[ 6162 ] = 8'h21;
  picture_data[ 6163 ] = 8'h01;
  picture_data[ 6164 ] = 8'h18;
  picture_data[ 6165 ] = 8'hE1;
  picture_data[ 6166 ] = 8'h21;
  picture_data[ 6167 ] = 8'h02;
  picture_data[ 6168 ] = 8'h20;
  picture_data[ 6169 ] = 8'hE2;
  picture_data[ 6170 ] = 8'h29;
  picture_data[ 6171 ] = 8'h02;
  picture_data[ 6172 ] = 8'h29;
  picture_data[ 6173 ] = 8'h23;
  picture_data[ 6174 ] = 8'h20;
  picture_data[ 6175 ] = 8'hE2;
  picture_data[ 6176 ] = 8'h21;
  picture_data[ 6177 ] = 8'h22;
  picture_data[ 6178 ] = 8'h31;
  picture_data[ 6179 ] = 8'hA4;
  picture_data[ 6180 ] = 8'h31;
  picture_data[ 6181 ] = 8'h83;
  picture_data[ 6182 ] = 8'h29;
  picture_data[ 6183 ] = 8'h62;
  picture_data[ 6184 ] = 8'h31;
  picture_data[ 6185 ] = 8'h83;
  picture_data[ 6186 ] = 8'h39;
  picture_data[ 6187 ] = 8'hA3;
  picture_data[ 6188 ] = 8'h29;
  picture_data[ 6189 ] = 8'h41;
  picture_data[ 6190 ] = 8'h39;
  picture_data[ 6191 ] = 8'hC3;
  picture_data[ 6192 ] = 8'h31;
  picture_data[ 6193 ] = 8'h82;
  picture_data[ 6194 ] = 8'h39;
  picture_data[ 6195 ] = 8'hA3;
  picture_data[ 6196 ] = 8'h29;
  picture_data[ 6197 ] = 8'h41;
  picture_data[ 6198 ] = 8'h31;
  picture_data[ 6199 ] = 8'h83;
  picture_data[ 6200 ] = 8'h29;
  picture_data[ 6201 ] = 8'h62;
  picture_data[ 6202 ] = 8'h31;
  picture_data[ 6203 ] = 8'h83;
  picture_data[ 6204 ] = 8'h39;
  picture_data[ 6205 ] = 8'hC4;
  picture_data[ 6206 ] = 8'h42;
  picture_data[ 6207 ] = 8'h25;
  picture_data[ 6208 ] = 8'h29;
  picture_data[ 6209 ] = 8'h62;
  picture_data[ 6210 ] = 8'h29;
  picture_data[ 6211 ] = 8'h42;
  picture_data[ 6212 ] = 8'h31;
  picture_data[ 6213 ] = 8'h83;
  picture_data[ 6214 ] = 8'h31;
  picture_data[ 6215 ] = 8'hA4;
  picture_data[ 6216 ] = 8'h42;
  picture_data[ 6217 ] = 8'h06;
  picture_data[ 6218 ] = 8'h29;
  picture_data[ 6219 ] = 8'h23;
  picture_data[ 6220 ] = 8'h29;
  picture_data[ 6221 ] = 8'h23;
  picture_data[ 6222 ] = 8'h20;
  picture_data[ 6223 ] = 8'hE2;
  picture_data[ 6224 ] = 8'h20;
  picture_data[ 6225 ] = 8'hE2;
  picture_data[ 6226 ] = 8'h29;
  picture_data[ 6227 ] = 8'h23;
  picture_data[ 6228 ] = 8'h29;
  picture_data[ 6229 ] = 8'h23;
  picture_data[ 6230 ] = 8'h08;
  picture_data[ 6231 ] = 8'hA8;
  picture_data[ 6232 ] = 8'h00;
  picture_data[ 6233 ] = 8'hA9;
  picture_data[ 6234 ] = 8'h00;
  picture_data[ 6235 ] = 8'hEF;
  picture_data[ 6236 ] = 8'h2A;
  picture_data[ 6237 ] = 8'hB8;
  picture_data[ 6238 ] = 8'h54;
  picture_data[ 6239 ] = 8'h3F;
  picture_data[ 6240 ] = 8'h22;
  picture_data[ 6241 ] = 8'h7A;
  picture_data[ 6242 ] = 8'h00;
  picture_data[ 6243 ] = 8'h90;
  picture_data[ 6244 ] = 8'h00;
  picture_data[ 6245 ] = 8'hCD;
  picture_data[ 6246 ] = 8'h19;
  picture_data[ 6247 ] = 8'h0A;
  picture_data[ 6248 ] = 8'h21;
  picture_data[ 6249 ] = 8'h28;
  picture_data[ 6250 ] = 8'h10;
  picture_data[ 6251 ] = 8'hE7;
  picture_data[ 6252 ] = 8'h10;
  picture_data[ 6253 ] = 8'hC7;
  picture_data[ 6254 ] = 8'h10;
  picture_data[ 6255 ] = 8'hC8;
  picture_data[ 6256 ] = 8'h10;
  picture_data[ 6257 ] = 8'hC7;
  picture_data[ 6258 ] = 8'h18;
  picture_data[ 6259 ] = 8'hC6;
  picture_data[ 6260 ] = 8'h08;
  picture_data[ 6261 ] = 8'h63;
  picture_data[ 6262 ] = 8'h10;
  picture_data[ 6263 ] = 8'hA3;
  picture_data[ 6264 ] = 8'h08;
  picture_data[ 6265 ] = 8'h81;
  picture_data[ 6266 ] = 8'h00;
  picture_data[ 6267 ] = 8'h20;
  picture_data[ 6268 ] = 8'h00;
  picture_data[ 6269 ] = 8'h20;
  picture_data[ 6270 ] = 8'h00;
  picture_data[ 6271 ] = 8'h61;
  picture_data[ 6272 ] = 8'h00;
  picture_data[ 6273 ] = 8'h60;
  picture_data[ 6274 ] = 8'h00;
  picture_data[ 6275 ] = 8'h60;
  picture_data[ 6276 ] = 8'h10;
  picture_data[ 6277 ] = 8'hC2;
  picture_data[ 6278 ] = 8'h10;
  picture_data[ 6279 ] = 8'hC2;
  picture_data[ 6280 ] = 8'h19;
  picture_data[ 6281 ] = 8'h03;
  picture_data[ 6282 ] = 8'h10;
  picture_data[ 6283 ] = 8'hC2;
  picture_data[ 6284 ] = 8'h08;
  picture_data[ 6285 ] = 8'h81;
  picture_data[ 6286 ] = 8'h10;
  picture_data[ 6287 ] = 8'hA1;
  picture_data[ 6288 ] = 8'h18;
  picture_data[ 6289 ] = 8'hC2;
  picture_data[ 6290 ] = 8'h18;
  picture_data[ 6291 ] = 8'hE2;
  picture_data[ 6292 ] = 8'h10;
  picture_data[ 6293 ] = 8'hA2;
  picture_data[ 6294 ] = 8'h18;
  picture_data[ 6295 ] = 8'hA1;
  picture_data[ 6296 ] = 8'h10;
  picture_data[ 6297 ] = 8'h80;
  picture_data[ 6298 ] = 8'h18;
  picture_data[ 6299 ] = 8'hA1;
  picture_data[ 6300 ] = 8'h18;
  picture_data[ 6301 ] = 8'hC1;
  picture_data[ 6302 ] = 8'h10;
  picture_data[ 6303 ] = 8'hA1;
  picture_data[ 6304 ] = 8'h18;
  picture_data[ 6305 ] = 8'hC1;
  picture_data[ 6306 ] = 8'h18;
  picture_data[ 6307 ] = 8'hC1;
  picture_data[ 6308 ] = 8'h18;
  picture_data[ 6309 ] = 8'hE2;
  picture_data[ 6310 ] = 8'h18;
  picture_data[ 6311 ] = 8'hC1;
  picture_data[ 6312 ] = 8'h18;
  picture_data[ 6313 ] = 8'hC1;
  picture_data[ 6314 ] = 8'h21;
  picture_data[ 6315 ] = 8'h02;
  picture_data[ 6316 ] = 8'h20;
  picture_data[ 6317 ] = 8'hE1;
  picture_data[ 6318 ] = 8'h29;
  picture_data[ 6319 ] = 8'h22;
  picture_data[ 6320 ] = 8'h20;
  picture_data[ 6321 ] = 8'hE2;
  picture_data[ 6322 ] = 8'h20;
  picture_data[ 6323 ] = 8'hC2;
  picture_data[ 6324 ] = 8'h29;
  picture_data[ 6325 ] = 8'h03;
  picture_data[ 6326 ] = 8'h31;
  picture_data[ 6327 ] = 8'h64;
  picture_data[ 6328 ] = 8'h42;
  picture_data[ 6329 ] = 8'h06;
  picture_data[ 6330 ] = 8'h29;
  picture_data[ 6331 ] = 8'h43;
  picture_data[ 6332 ] = 8'h18;
  picture_data[ 6333 ] = 8'hC0;
  picture_data[ 6334 ] = 8'h29;
  picture_data[ 6335 ] = 8'h42;
  picture_data[ 6336 ] = 8'h31;
  picture_data[ 6337 ] = 8'h63;
  picture_data[ 6338 ] = 8'h31;
  picture_data[ 6339 ] = 8'h62;
  picture_data[ 6340 ] = 8'h31;
  picture_data[ 6341 ] = 8'h82;
  picture_data[ 6342 ] = 8'h39;
  picture_data[ 6343 ] = 8'hA3;
  picture_data[ 6344 ] = 8'h31;
  picture_data[ 6345 ] = 8'h82;
  picture_data[ 6346 ] = 8'h31;
  picture_data[ 6347 ] = 8'h82;
  picture_data[ 6348 ] = 8'h31;
  picture_data[ 6349 ] = 8'h62;
  picture_data[ 6350 ] = 8'h42;
  picture_data[ 6351 ] = 8'h04;
  picture_data[ 6352 ] = 8'h29;
  picture_data[ 6353 ] = 8'h41;
  picture_data[ 6354 ] = 8'h42;
  picture_data[ 6355 ] = 8'h05;
  picture_data[ 6356 ] = 8'h5A;
  picture_data[ 6357 ] = 8'hA7;
  picture_data[ 6358 ] = 8'h42;
  picture_data[ 6359 ] = 8'h25;
  picture_data[ 6360 ] = 8'h42;
  picture_data[ 6361 ] = 8'h45;
  picture_data[ 6362 ] = 8'h39;
  picture_data[ 6363 ] = 8'hC4;
  picture_data[ 6364 ] = 8'h29;
  picture_data[ 6365 ] = 8'h83;
  picture_data[ 6366 ] = 8'h31;
  picture_data[ 6367 ] = 8'hA4;
  picture_data[ 6368 ] = 8'h21;
  picture_data[ 6369 ] = 8'h23;
  picture_data[ 6370 ] = 8'h29;
  picture_data[ 6371 ] = 8'h43;
  picture_data[ 6372 ] = 8'h29;
  picture_data[ 6373 ] = 8'h23;
  picture_data[ 6374 ] = 8'h10;
  picture_data[ 6375 ] = 8'hA1;
  picture_data[ 6376 ] = 8'h10;
  picture_data[ 6377 ] = 8'h81;
  picture_data[ 6378 ] = 8'h18;
  picture_data[ 6379 ] = 8'hC2;
  picture_data[ 6380 ] = 8'h21;
  picture_data[ 6381 ] = 8'h02;
  picture_data[ 6382 ] = 8'h08;
  picture_data[ 6383 ] = 8'hA6;
  picture_data[ 6384 ] = 8'h00;
  picture_data[ 6385 ] = 8'h46;
  picture_data[ 6386 ] = 8'h00;
  picture_data[ 6387 ] = 8'hAA;
  picture_data[ 6388 ] = 8'h00;
  picture_data[ 6389 ] = 8'hCD;
  picture_data[ 6390 ] = 8'h01;
  picture_data[ 6391 ] = 8'h0F;
  picture_data[ 6392 ] = 8'h00;
  picture_data[ 6393 ] = 8'hAE;
  picture_data[ 6394 ] = 8'h00;
  picture_data[ 6395 ] = 8'h6C;
  picture_data[ 6396 ] = 8'h08;
  picture_data[ 6397 ] = 8'hCB;
  picture_data[ 6398 ] = 8'h00;
  picture_data[ 6399 ] = 8'h86;
  picture_data[ 6400 ] = 8'h00;
  picture_data[ 6401 ] = 8'h65;
  picture_data[ 6402 ] = 8'h10;
  picture_data[ 6403 ] = 8'hA7;
  picture_data[ 6404 ] = 8'h19;
  picture_data[ 6405 ] = 8'h09;
  picture_data[ 6406 ] = 8'h19;
  picture_data[ 6407 ] = 8'h0A;
  picture_data[ 6408 ] = 8'h21;
  picture_data[ 6409 ] = 8'h2A;
  picture_data[ 6410 ] = 8'h18;
  picture_data[ 6411 ] = 8'hC8;
  picture_data[ 6412 ] = 8'h08;
  picture_data[ 6413 ] = 8'h65;
  picture_data[ 6414 ] = 8'h08;
  picture_data[ 6415 ] = 8'h83;
  picture_data[ 6416 ] = 8'h08;
  picture_data[ 6417 ] = 8'h81;
  picture_data[ 6418 ] = 8'h00;
  picture_data[ 6419 ] = 8'h41;
  picture_data[ 6420 ] = 8'h00;
  picture_data[ 6421 ] = 8'h61;
  picture_data[ 6422 ] = 8'h00;
  picture_data[ 6423 ] = 8'h61;
  picture_data[ 6424 ] = 8'h00;
  picture_data[ 6425 ] = 8'h41;
  picture_data[ 6426 ] = 8'h00;
  picture_data[ 6427 ] = 8'h81;
  picture_data[ 6428 ] = 8'h10;
  picture_data[ 6429 ] = 8'hE3;
  picture_data[ 6430 ] = 8'h10;
  picture_data[ 6431 ] = 8'hA2;
  picture_data[ 6432 ] = 8'h10;
  picture_data[ 6433 ] = 8'hA2;
  picture_data[ 6434 ] = 8'h08;
  picture_data[ 6435 ] = 8'h81;
  picture_data[ 6436 ] = 8'h08;
  picture_data[ 6437 ] = 8'hA1;
  picture_data[ 6438 ] = 8'h10;
  picture_data[ 6439 ] = 8'h81;
  picture_data[ 6440 ] = 8'h08;
  picture_data[ 6441 ] = 8'h40;
  picture_data[ 6442 ] = 8'h10;
  picture_data[ 6443 ] = 8'h61;
  picture_data[ 6444 ] = 8'h18;
  picture_data[ 6445 ] = 8'hC2;
  picture_data[ 6446 ] = 8'h10;
  picture_data[ 6447 ] = 8'hC2;
  picture_data[ 6448 ] = 8'h10;
  picture_data[ 6449 ] = 8'hA1;
  picture_data[ 6450 ] = 8'h10;
  picture_data[ 6451 ] = 8'hC1;
  picture_data[ 6452 ] = 8'h10;
  picture_data[ 6453 ] = 8'hC0;
  picture_data[ 6454 ] = 8'h18;
  picture_data[ 6455 ] = 8'hE1;
  picture_data[ 6456 ] = 8'h19;
  picture_data[ 6457 ] = 8'h01;
  picture_data[ 6458 ] = 8'h18;
  picture_data[ 6459 ] = 8'hE1;
  picture_data[ 6460 ] = 8'h19;
  picture_data[ 6461 ] = 8'h02;
  picture_data[ 6462 ] = 8'h21;
  picture_data[ 6463 ] = 8'h22;
  picture_data[ 6464 ] = 8'h18;
  picture_data[ 6465 ] = 8'hE1;
  picture_data[ 6466 ] = 8'h18;
  picture_data[ 6467 ] = 8'hC0;
  picture_data[ 6468 ] = 8'h20;
  picture_data[ 6469 ] = 8'hE1;
  picture_data[ 6470 ] = 8'h18;
  picture_data[ 6471 ] = 8'hE1;
  picture_data[ 6472 ] = 8'h18;
  picture_data[ 6473 ] = 8'hC0;
  picture_data[ 6474 ] = 8'h21;
  picture_data[ 6475 ] = 8'h23;
  picture_data[ 6476 ] = 8'h20;
  picture_data[ 6477 ] = 8'hE2;
  picture_data[ 6478 ] = 8'h29;
  picture_data[ 6479 ] = 8'h02;
  picture_data[ 6480 ] = 8'h39;
  picture_data[ 6481 ] = 8'hA4;
  picture_data[ 6482 ] = 8'h29;
  picture_data[ 6483 ] = 8'h22;
  picture_data[ 6484 ] = 8'h18;
  picture_data[ 6485 ] = 8'hA0;
  picture_data[ 6486 ] = 8'h39;
  picture_data[ 6487 ] = 8'h83;
  picture_data[ 6488 ] = 8'h29;
  picture_data[ 6489 ] = 8'h42;
  picture_data[ 6490 ] = 8'h39;
  picture_data[ 6491 ] = 8'hC3;
  picture_data[ 6492 ] = 8'h41;
  picture_data[ 6493 ] = 8'hE4;
  picture_data[ 6494 ] = 8'h31;
  picture_data[ 6495 ] = 8'h62;
  picture_data[ 6496 ] = 8'h31;
  picture_data[ 6497 ] = 8'h62;
  picture_data[ 6498 ] = 8'h31;
  picture_data[ 6499 ] = 8'h82;
  picture_data[ 6500 ] = 8'h31;
  picture_data[ 6501 ] = 8'h82;
  picture_data[ 6502 ] = 8'h41;
  picture_data[ 6503 ] = 8'hE4;
  picture_data[ 6504 ] = 8'h39;
  picture_data[ 6505 ] = 8'h83;
  picture_data[ 6506 ] = 8'h31;
  picture_data[ 6507 ] = 8'h82;
  picture_data[ 6508 ] = 8'h52;
  picture_data[ 6509 ] = 8'h86;
  picture_data[ 6510 ] = 8'h4A;
  picture_data[ 6511 ] = 8'h66;
  picture_data[ 6512 ] = 8'h3A;
  picture_data[ 6513 ] = 8'h04;
  picture_data[ 6514 ] = 8'h42;
  picture_data[ 6515 ] = 8'h26;
  picture_data[ 6516 ] = 8'h39;
  picture_data[ 6517 ] = 8'hE4;
  picture_data[ 6518 ] = 8'h29;
  picture_data[ 6519 ] = 8'h84;
  picture_data[ 6520 ] = 8'h19;
  picture_data[ 6521 ] = 8'h02;
  picture_data[ 6522 ] = 8'h29;
  picture_data[ 6523 ] = 8'h43;
  picture_data[ 6524 ] = 8'h21;
  picture_data[ 6525 ] = 8'h23;
  picture_data[ 6526 ] = 8'h21;
  picture_data[ 6527 ] = 8'h02;
  picture_data[ 6528 ] = 8'h18;
  picture_data[ 6529 ] = 8'hC1;
  picture_data[ 6530 ] = 8'h18;
  picture_data[ 6531 ] = 8'hC1;
  picture_data[ 6532 ] = 8'h10;
  picture_data[ 6533 ] = 8'hA1;
  picture_data[ 6534 ] = 8'h08;
  picture_data[ 6535 ] = 8'h85;
  picture_data[ 6536 ] = 8'h10;
  picture_data[ 6537 ] = 8'hE8;
  picture_data[ 6538 ] = 8'h08;
  picture_data[ 6539 ] = 8'hA8;
  picture_data[ 6540 ] = 8'h08;
  picture_data[ 6541 ] = 8'hCA;
  picture_data[ 6542 ] = 8'h00;
  picture_data[ 6543 ] = 8'h8A;
  picture_data[ 6544 ] = 8'h00;
  picture_data[ 6545 ] = 8'hAA;
  picture_data[ 6546 ] = 8'h11;
  picture_data[ 6547 ] = 8'h0B;
  picture_data[ 6548 ] = 8'h10;
  picture_data[ 6549 ] = 8'hEA;
  picture_data[ 6550 ] = 8'h19;
  picture_data[ 6551 ] = 8'h29;
  picture_data[ 6552 ] = 8'h10;
  picture_data[ 6553 ] = 8'hE7;
  picture_data[ 6554 ] = 8'h08;
  picture_data[ 6555 ] = 8'h86;
  picture_data[ 6556 ] = 8'h08;
  picture_data[ 6557 ] = 8'hA7;
  picture_data[ 6558 ] = 8'h10;
  picture_data[ 6559 ] = 8'hA8;
  picture_data[ 6560 ] = 8'h08;
  picture_data[ 6561 ] = 8'h87;
  picture_data[ 6562 ] = 8'h29;
  picture_data[ 6563 ] = 8'h6B;
  picture_data[ 6564 ] = 8'h10;
  picture_data[ 6565 ] = 8'hA6;
  picture_data[ 6566 ] = 8'h00;
  picture_data[ 6567 ] = 8'h63;
  picture_data[ 6568 ] = 8'h00;
  picture_data[ 6569 ] = 8'h61;
  picture_data[ 6570 ] = 8'h00;
  picture_data[ 6571 ] = 8'h61;
  picture_data[ 6572 ] = 8'h00;
  picture_data[ 6573 ] = 8'h81;
  picture_data[ 6574 ] = 8'h08;
  picture_data[ 6575 ] = 8'h82;
  picture_data[ 6576 ] = 8'h00;
  picture_data[ 6577 ] = 8'h61;
  picture_data[ 6578 ] = 8'h00;
  picture_data[ 6579 ] = 8'h61;
  picture_data[ 6580 ] = 8'h10;
  picture_data[ 6581 ] = 8'hA2;
  picture_data[ 6582 ] = 8'h08;
  picture_data[ 6583 ] = 8'h61;
  picture_data[ 6584 ] = 8'h10;
  picture_data[ 6585 ] = 8'hA2;
  picture_data[ 6586 ] = 8'h10;
  picture_data[ 6587 ] = 8'hC2;
  picture_data[ 6588 ] = 8'h10;
  picture_data[ 6589 ] = 8'hC2;
  picture_data[ 6590 ] = 8'h10;
  picture_data[ 6591 ] = 8'hA2;
  picture_data[ 6592 ] = 8'h08;
  picture_data[ 6593 ] = 8'h61;
  picture_data[ 6594 ] = 8'h10;
  picture_data[ 6595 ] = 8'h81;
  picture_data[ 6596 ] = 8'h10;
  picture_data[ 6597 ] = 8'hA2;
  picture_data[ 6598 ] = 8'h10;
  picture_data[ 6599 ] = 8'hC2;
  picture_data[ 6600 ] = 8'h19;
  picture_data[ 6601 ] = 8'h03;
  picture_data[ 6602 ] = 8'h10;
  picture_data[ 6603 ] = 8'hC1;
  picture_data[ 6604 ] = 8'h08;
  picture_data[ 6605 ] = 8'h80;
  picture_data[ 6606 ] = 8'h10;
  picture_data[ 6607 ] = 8'hC0;
  picture_data[ 6608 ] = 8'h19;
  picture_data[ 6609 ] = 8'h02;
  picture_data[ 6610 ] = 8'h18;
  picture_data[ 6611 ] = 8'hE2;
  picture_data[ 6612 ] = 8'h18;
  picture_data[ 6613 ] = 8'hE1;
  picture_data[ 6614 ] = 8'h21;
  picture_data[ 6615 ] = 8'h02;
  picture_data[ 6616 ] = 8'h10;
  picture_data[ 6617 ] = 8'hA0;
  picture_data[ 6618 ] = 8'h18;
  picture_data[ 6619 ] = 8'hC0;
  picture_data[ 6620 ] = 8'h10;
  picture_data[ 6621 ] = 8'hA0;
  picture_data[ 6622 ] = 8'h10;
  picture_data[ 6623 ] = 8'hA0;
  picture_data[ 6624 ] = 8'h21;
  picture_data[ 6625 ] = 8'h02;
  picture_data[ 6626 ] = 8'h29;
  picture_data[ 6627 ] = 8'h43;
  picture_data[ 6628 ] = 8'h31;
  picture_data[ 6629 ] = 8'h43;
  picture_data[ 6630 ] = 8'h18;
  picture_data[ 6631 ] = 8'h80;
  picture_data[ 6632 ] = 8'h20;
  picture_data[ 6633 ] = 8'hA0;
  picture_data[ 6634 ] = 8'h39;
  picture_data[ 6635 ] = 8'h83;
  picture_data[ 6636 ] = 8'h39;
  picture_data[ 6637 ] = 8'h83;
  picture_data[ 6638 ] = 8'h20;
  picture_data[ 6639 ] = 8'hE0;
  picture_data[ 6640 ] = 8'h20;
  picture_data[ 6641 ] = 8'hE0;
  picture_data[ 6642 ] = 8'h52;
  picture_data[ 6643 ] = 8'h46;
  picture_data[ 6644 ] = 8'h4A;
  picture_data[ 6645 ] = 8'h45;
  picture_data[ 6646 ] = 8'h29;
  picture_data[ 6647 ] = 8'h21;
  picture_data[ 6648 ] = 8'h39;
  picture_data[ 6649 ] = 8'hA3;
  picture_data[ 6650 ] = 8'h31;
  picture_data[ 6651 ] = 8'h83;
  picture_data[ 6652 ] = 8'h31;
  picture_data[ 6653 ] = 8'h62;
  picture_data[ 6654 ] = 8'h41;
  picture_data[ 6655 ] = 8'hC4;
  picture_data[ 6656 ] = 8'h42;
  picture_data[ 6657 ] = 8'h04;
  picture_data[ 6658 ] = 8'h31;
  picture_data[ 6659 ] = 8'h42;
  picture_data[ 6660 ] = 8'h31;
  picture_data[ 6661 ] = 8'h62;
  picture_data[ 6662 ] = 8'h4A;
  picture_data[ 6663 ] = 8'h66;
  picture_data[ 6664 ] = 8'h3A;
  picture_data[ 6665 ] = 8'h05;
  picture_data[ 6666 ] = 8'h3A;
  picture_data[ 6667 ] = 8'h05;
  picture_data[ 6668 ] = 8'h31;
  picture_data[ 6669 ] = 8'hC4;
  picture_data[ 6670 ] = 8'h21;
  picture_data[ 6671 ] = 8'h22;
  picture_data[ 6672 ] = 8'h19;
  picture_data[ 6673 ] = 8'h02;
  picture_data[ 6674 ] = 8'h19;
  picture_data[ 6675 ] = 8'h02;
  picture_data[ 6676 ] = 8'h18;
  picture_data[ 6677 ] = 8'hE2;
  picture_data[ 6678 ] = 8'h19;
  picture_data[ 6679 ] = 8'h02;
  picture_data[ 6680 ] = 8'h18;
  picture_data[ 6681 ] = 8'hE1;
  picture_data[ 6682 ] = 8'h21;
  picture_data[ 6683 ] = 8'h22;
  picture_data[ 6684 ] = 8'h21;
  picture_data[ 6685 ] = 8'h42;
  picture_data[ 6686 ] = 8'h00;
  picture_data[ 6687 ] = 8'h45;
  picture_data[ 6688 ] = 8'h08;
  picture_data[ 6689 ] = 8'h85;
  picture_data[ 6690 ] = 8'h00;
  picture_data[ 6691 ] = 8'h25;
  picture_data[ 6692 ] = 8'h08;
  picture_data[ 6693 ] = 8'hA7;
  picture_data[ 6694 ] = 8'h10;
  picture_data[ 6695 ] = 8'hE8;
  picture_data[ 6696 ] = 8'h10;
  picture_data[ 6697 ] = 8'hC8;
  picture_data[ 6698 ] = 8'h08;
  picture_data[ 6699 ] = 8'hA8;
  picture_data[ 6700 ] = 8'h19;
  picture_data[ 6701 ] = 8'h09;
  picture_data[ 6702 ] = 8'h19;
  picture_data[ 6703 ] = 8'h48;
  picture_data[ 6704 ] = 8'h10;
  picture_data[ 6705 ] = 8'hE6;
  picture_data[ 6706 ] = 8'h19;
  picture_data[ 6707 ] = 8'h27;
  picture_data[ 6708 ] = 8'h08;
  picture_data[ 6709 ] = 8'hA5;
  picture_data[ 6710 ] = 8'h08;
  picture_data[ 6711 ] = 8'h84;
  picture_data[ 6712 ] = 8'h08;
  picture_data[ 6713 ] = 8'hA4;
  picture_data[ 6714 ] = 8'h19;
  picture_data[ 6715 ] = 8'h06;
  picture_data[ 6716 ] = 8'h08;
  picture_data[ 6717 ] = 8'h84;
  picture_data[ 6718 ] = 8'h08;
  picture_data[ 6719 ] = 8'hA3;
  picture_data[ 6720 ] = 8'h08;
  picture_data[ 6721 ] = 8'h82;
  picture_data[ 6722 ] = 8'h00;
  picture_data[ 6723 ] = 8'h61;
  picture_data[ 6724 ] = 8'h00;
  picture_data[ 6725 ] = 8'h41;
  picture_data[ 6726 ] = 8'h08;
  picture_data[ 6727 ] = 8'h61;
  picture_data[ 6728 ] = 8'h08;
  picture_data[ 6729 ] = 8'h61;
  picture_data[ 6730 ] = 8'h00;
  picture_data[ 6731 ] = 8'h61;
  picture_data[ 6732 ] = 8'h00;
  picture_data[ 6733 ] = 8'h41;
  picture_data[ 6734 ] = 8'h00;
  picture_data[ 6735 ] = 8'h61;
  picture_data[ 6736 ] = 8'h08;
  picture_data[ 6737 ] = 8'h81;
  picture_data[ 6738 ] = 8'h08;
  picture_data[ 6739 ] = 8'hA1;
  picture_data[ 6740 ] = 8'h18;
  picture_data[ 6741 ] = 8'hE3;
  picture_data[ 6742 ] = 8'h18;
  picture_data[ 6743 ] = 8'hE3;
  picture_data[ 6744 ] = 8'h10;
  picture_data[ 6745 ] = 8'h81;
  picture_data[ 6746 ] = 8'h08;
  picture_data[ 6747 ] = 8'h40;
  picture_data[ 6748 ] = 8'h00;
  picture_data[ 6749 ] = 8'h40;
  picture_data[ 6750 ] = 8'h08;
  picture_data[ 6751 ] = 8'h81;
  picture_data[ 6752 ] = 8'h18;
  picture_data[ 6753 ] = 8'hE2;
  picture_data[ 6754 ] = 8'h10;
  picture_data[ 6755 ] = 8'hC1;
  picture_data[ 6756 ] = 8'h08;
  picture_data[ 6757 ] = 8'h80;
  picture_data[ 6758 ] = 8'h10;
  picture_data[ 6759 ] = 8'hC1;
  picture_data[ 6760 ] = 8'h19;
  picture_data[ 6761 ] = 8'h03;
  picture_data[ 6762 ] = 8'h21;
  picture_data[ 6763 ] = 8'h03;
  picture_data[ 6764 ] = 8'h20;
  picture_data[ 6765 ] = 8'hE3;
  picture_data[ 6766 ] = 8'h18;
  picture_data[ 6767 ] = 8'hA2;
  picture_data[ 6768 ] = 8'h18;
  picture_data[ 6769 ] = 8'hC2;
  picture_data[ 6770 ] = 8'h18;
  picture_data[ 6771 ] = 8'hA1;
  picture_data[ 6772 ] = 8'h18;
  picture_data[ 6773 ] = 8'hA1;
  picture_data[ 6774 ] = 8'h18;
  picture_data[ 6775 ] = 8'hC0;
  picture_data[ 6776 ] = 8'h29;
  picture_data[ 6777 ] = 8'h22;
  picture_data[ 6778 ] = 8'h31;
  picture_data[ 6779 ] = 8'h63;
  picture_data[ 6780 ] = 8'h31;
  picture_data[ 6781 ] = 8'h21;
  picture_data[ 6782 ] = 8'h30;
  picture_data[ 6783 ] = 8'hE0;
  picture_data[ 6784 ] = 8'h49;
  picture_data[ 6785 ] = 8'h82;
  picture_data[ 6786 ] = 8'h49;
  picture_data[ 6787 ] = 8'hA3;
  picture_data[ 6788 ] = 8'h41;
  picture_data[ 6789 ] = 8'h83;
  picture_data[ 6790 ] = 8'h31;
  picture_data[ 6791 ] = 8'h00;
  picture_data[ 6792 ] = 8'h39;
  picture_data[ 6793 ] = 8'h62;
  picture_data[ 6794 ] = 8'h31;
  picture_data[ 6795 ] = 8'h82;
  picture_data[ 6796 ] = 8'h39;
  picture_data[ 6797 ] = 8'hA3;
  picture_data[ 6798 ] = 8'h29;
  picture_data[ 6799 ] = 8'h42;
  picture_data[ 6800 ] = 8'h41;
  picture_data[ 6801 ] = 8'hE4;
  picture_data[ 6802 ] = 8'h39;
  picture_data[ 6803 ] = 8'hC4;
  picture_data[ 6804 ] = 8'h29;
  picture_data[ 6805 ] = 8'h42;
  picture_data[ 6806 ] = 8'h42;
  picture_data[ 6807 ] = 8'h05;
  picture_data[ 6808 ] = 8'h52;
  picture_data[ 6809 ] = 8'h87;
  picture_data[ 6810 ] = 8'h41;
  picture_data[ 6811 ] = 8'hE4;
  picture_data[ 6812 ] = 8'h29;
  picture_data[ 6813 ] = 8'h41;
  picture_data[ 6814 ] = 8'h31;
  picture_data[ 6815 ] = 8'h83;
  picture_data[ 6816 ] = 8'h52;
  picture_data[ 6817 ] = 8'h87;
  picture_data[ 6818 ] = 8'h31;
  picture_data[ 6819 ] = 8'hA4;
  picture_data[ 6820 ] = 8'h21;
  picture_data[ 6821 ] = 8'h43;
  picture_data[ 6822 ] = 8'h19;
  picture_data[ 6823 ] = 8'h02;
  picture_data[ 6824 ] = 8'h18;
  picture_data[ 6825 ] = 8'hE2;
  picture_data[ 6826 ] = 8'h19;
  picture_data[ 6827 ] = 8'h02;
  picture_data[ 6828 ] = 8'h21;
  picture_data[ 6829 ] = 8'h22;
  picture_data[ 6830 ] = 8'h21;
  picture_data[ 6831 ] = 8'h63;
  picture_data[ 6832 ] = 8'h21;
  picture_data[ 6833 ] = 8'h22;
  picture_data[ 6834 ] = 8'h21;
  picture_data[ 6835 ] = 8'h43;
  picture_data[ 6836 ] = 8'h21;
  picture_data[ 6837 ] = 8'h63;
  picture_data[ 6838 ] = 8'h08;
  picture_data[ 6839 ] = 8'h85;
  picture_data[ 6840 ] = 8'h00;
  picture_data[ 6841 ] = 8'h44;
  picture_data[ 6842 ] = 8'h18;
  picture_data[ 6843 ] = 8'hE6;
  picture_data[ 6844 ] = 8'h10;
  picture_data[ 6845 ] = 8'hC6;
  picture_data[ 6846 ] = 8'h21;
  picture_data[ 6847 ] = 8'h48;
  picture_data[ 6848 ] = 8'h29;
  picture_data[ 6849 ] = 8'h69;
  picture_data[ 6850 ] = 8'h19;
  picture_data[ 6851 ] = 8'h09;
  picture_data[ 6852 ] = 8'h19;
  picture_data[ 6853 ] = 8'h09;
  picture_data[ 6854 ] = 8'h10;
  picture_data[ 6855 ] = 8'hC6;
  picture_data[ 6856 ] = 8'h08;
  picture_data[ 6857 ] = 8'hA5;
  picture_data[ 6858 ] = 8'h00;
  picture_data[ 6859 ] = 8'h63;
  picture_data[ 6860 ] = 8'h08;
  picture_data[ 6861 ] = 8'hA4;
  picture_data[ 6862 ] = 8'h00;
  picture_data[ 6863 ] = 8'h62;
  picture_data[ 6864 ] = 8'h00;
  picture_data[ 6865 ] = 8'h21;
  picture_data[ 6866 ] = 8'h08;
  picture_data[ 6867 ] = 8'hC3;
  picture_data[ 6868 ] = 8'h08;
  picture_data[ 6869 ] = 8'h83;
  picture_data[ 6870 ] = 8'h08;
  picture_data[ 6871 ] = 8'hA3;
  picture_data[ 6872 ] = 8'h10;
  picture_data[ 6873 ] = 8'hA3;
  picture_data[ 6874 ] = 8'h10;
  picture_data[ 6875 ] = 8'hA2;
  picture_data[ 6876 ] = 8'h08;
  picture_data[ 6877 ] = 8'h62;
  picture_data[ 6878 ] = 8'h00;
  picture_data[ 6879 ] = 8'h41;
  picture_data[ 6880 ] = 8'h00;
  picture_data[ 6881 ] = 8'h41;
  picture_data[ 6882 ] = 8'h08;
  picture_data[ 6883 ] = 8'h61;
  picture_data[ 6884 ] = 8'h08;
  picture_data[ 6885 ] = 8'h61;
  picture_data[ 6886 ] = 8'h08;
  picture_data[ 6887 ] = 8'hA2;
  picture_data[ 6888 ] = 8'h08;
  picture_data[ 6889 ] = 8'h81;
  picture_data[ 6890 ] = 8'h08;
  picture_data[ 6891 ] = 8'hA1;
  picture_data[ 6892 ] = 8'h19;
  picture_data[ 6893 ] = 8'h03;
  picture_data[ 6894 ] = 8'h19;
  picture_data[ 6895 ] = 8'h03;
  picture_data[ 6896 ] = 8'h08;
  picture_data[ 6897 ] = 8'h61;
  picture_data[ 6898 ] = 8'h00;
  picture_data[ 6899 ] = 8'h40;
  picture_data[ 6900 ] = 8'h08;
  picture_data[ 6901 ] = 8'h60;
  picture_data[ 6902 ] = 8'h08;
  picture_data[ 6903 ] = 8'h60;
  picture_data[ 6904 ] = 8'h10;
  picture_data[ 6905 ] = 8'hC2;
  picture_data[ 6906 ] = 8'h08;
  picture_data[ 6907 ] = 8'hA1;
  picture_data[ 6908 ] = 8'h08;
  picture_data[ 6909 ] = 8'hA1;
  picture_data[ 6910 ] = 8'h10;
  picture_data[ 6911 ] = 8'hE2;
  picture_data[ 6912 ] = 8'h18;
  picture_data[ 6913 ] = 8'hE2;
  picture_data[ 6914 ] = 8'h18;
  picture_data[ 6915 ] = 8'hE3;
  picture_data[ 6916 ] = 8'h21;
  picture_data[ 6917 ] = 8'h03;
  picture_data[ 6918 ] = 8'h18;
  picture_data[ 6919 ] = 8'hA2;
  picture_data[ 6920 ] = 8'h31;
  picture_data[ 6921 ] = 8'h44;
  picture_data[ 6922 ] = 8'h18;
  picture_data[ 6923 ] = 8'hC1;
  picture_data[ 6924 ] = 8'h18;
  picture_data[ 6925 ] = 8'hA0;
  picture_data[ 6926 ] = 8'h29;
  picture_data[ 6927 ] = 8'h22;
  picture_data[ 6928 ] = 8'h29;
  picture_data[ 6929 ] = 8'h21;
  picture_data[ 6930 ] = 8'h28;
  picture_data[ 6931 ] = 8'hC0;
  picture_data[ 6932 ] = 8'h39;
  picture_data[ 6933 ] = 8'h21;
  picture_data[ 6934 ] = 8'h51;
  picture_data[ 6935 ] = 8'hA2;
  picture_data[ 6936 ] = 8'h41;
  picture_data[ 6937 ] = 8'h20;
  picture_data[ 6938 ] = 8'h49;
  picture_data[ 6939 ] = 8'h62;
  picture_data[ 6940 ] = 8'h41;
  picture_data[ 6941 ] = 8'h62;
  picture_data[ 6942 ] = 8'h39;
  picture_data[ 6943 ] = 8'h21;
  picture_data[ 6944 ] = 8'h39;
  picture_data[ 6945 ] = 8'h42;
  picture_data[ 6946 ] = 8'h41;
  picture_data[ 6947 ] = 8'hA3;
  picture_data[ 6948 ] = 8'h39;
  picture_data[ 6949 ] = 8'hA3;
  picture_data[ 6950 ] = 8'h39;
  picture_data[ 6951 ] = 8'hA3;
  picture_data[ 6952 ] = 8'h39;
  picture_data[ 6953 ] = 8'hC4;
  picture_data[ 6954 ] = 8'h4A;
  picture_data[ 6955 ] = 8'h05;
  picture_data[ 6956 ] = 8'h39;
  picture_data[ 6957 ] = 8'hA4;
  picture_data[ 6958 ] = 8'h39;
  picture_data[ 6959 ] = 8'h83;
  picture_data[ 6960 ] = 8'h6B;
  picture_data[ 6961 ] = 8'h09;
  picture_data[ 6962 ] = 8'h39;
  picture_data[ 6963 ] = 8'hA3;
  picture_data[ 6964 ] = 8'h31;
  picture_data[ 6965 ] = 8'h83;
  picture_data[ 6966 ] = 8'h20;
  picture_data[ 6967 ] = 8'hC1;
  picture_data[ 6968 ] = 8'h39;
  picture_data[ 6969 ] = 8'hA4;
  picture_data[ 6970 ] = 8'h29;
  picture_data[ 6971 ] = 8'h43;
  picture_data[ 6972 ] = 8'h18;
  picture_data[ 6973 ] = 8'hE2;
  picture_data[ 6974 ] = 8'h20;
  picture_data[ 6975 ] = 8'hE2;
  picture_data[ 6976 ] = 8'h21;
  picture_data[ 6977 ] = 8'h02;
  picture_data[ 6978 ] = 8'h19;
  picture_data[ 6979 ] = 8'h02;
  picture_data[ 6980 ] = 8'h21;
  picture_data[ 6981 ] = 8'h23;
  picture_data[ 6982 ] = 8'h21;
  picture_data[ 6983 ] = 8'h23;
  picture_data[ 6984 ] = 8'h19;
  picture_data[ 6985 ] = 8'h01;
  picture_data[ 6986 ] = 8'h18;
  picture_data[ 6987 ] = 8'hE1;
  picture_data[ 6988 ] = 8'h18;
  picture_data[ 6989 ] = 8'hE1;
  picture_data[ 6990 ] = 8'h10;
  picture_data[ 6991 ] = 8'hA5;
  picture_data[ 6992 ] = 8'h10;
  picture_data[ 6993 ] = 8'hE5;
  picture_data[ 6994 ] = 8'h10;
  picture_data[ 6995 ] = 8'hE5;
  picture_data[ 6996 ] = 8'h19;
  picture_data[ 6997 ] = 8'h46;
  picture_data[ 6998 ] = 8'h29;
  picture_data[ 6999 ] = 8'hC9;
  picture_data[ 7000 ] = 8'h21;
  picture_data[ 7001 ] = 8'h69;
  picture_data[ 7002 ] = 8'h21;
  picture_data[ 7003 ] = 8'h4B;
  picture_data[ 7004 ] = 8'h18;
  picture_data[ 7005 ] = 8'hEA;
  picture_data[ 7006 ] = 8'h10;
  picture_data[ 7007 ] = 8'hC8;
  picture_data[ 7008 ] = 8'h08;
  picture_data[ 7009 ] = 8'h65;
  picture_data[ 7010 ] = 8'h08;
  picture_data[ 7011 ] = 8'h85;
  picture_data[ 7012 ] = 8'h08;
  picture_data[ 7013 ] = 8'hA5;
  picture_data[ 7014 ] = 8'h08;
  picture_data[ 7015 ] = 8'hA3;
  picture_data[ 7016 ] = 8'h00;
  picture_data[ 7017 ] = 8'h82;
  picture_data[ 7018 ] = 8'h00;
  picture_data[ 7019 ] = 8'h62;
  picture_data[ 7020 ] = 8'h08;
  picture_data[ 7021 ] = 8'hC3;
  picture_data[ 7022 ] = 8'h08;
  picture_data[ 7023 ] = 8'h62;
  picture_data[ 7024 ] = 8'h08;
  picture_data[ 7025 ] = 8'h62;
  picture_data[ 7026 ] = 8'h10;
  picture_data[ 7027 ] = 8'h82;
  picture_data[ 7028 ] = 8'h08;
  picture_data[ 7029 ] = 8'h62;
  picture_data[ 7030 ] = 8'h00;
  picture_data[ 7031 ] = 8'h41;
  picture_data[ 7032 ] = 8'h00;
  picture_data[ 7033 ] = 8'h20;
  picture_data[ 7034 ] = 8'h00;
  picture_data[ 7035 ] = 8'h40;
  picture_data[ 7036 ] = 8'h08;
  picture_data[ 7037 ] = 8'h41;
  picture_data[ 7038 ] = 8'h00;
  picture_data[ 7039 ] = 8'h40;
  picture_data[ 7040 ] = 8'h10;
  picture_data[ 7041 ] = 8'hA2;
  picture_data[ 7042 ] = 8'h10;
  picture_data[ 7043 ] = 8'hA2;
  picture_data[ 7044 ] = 8'h08;
  picture_data[ 7045 ] = 8'hA1;
  picture_data[ 7046 ] = 8'h08;
  picture_data[ 7047 ] = 8'h81;
  picture_data[ 7048 ] = 8'h08;
  picture_data[ 7049 ] = 8'hA1;
  picture_data[ 7050 ] = 8'h08;
  picture_data[ 7051 ] = 8'h80;
  picture_data[ 7052 ] = 8'h00;
  picture_data[ 7053 ] = 8'h40;
  picture_data[ 7054 ] = 8'h08;
  picture_data[ 7055 ] = 8'h61;
  picture_data[ 7056 ] = 8'h10;
  picture_data[ 7057 ] = 8'hC2;
  picture_data[ 7058 ] = 8'h08;
  picture_data[ 7059 ] = 8'hC2;
  picture_data[ 7060 ] = 8'h08;
  picture_data[ 7061 ] = 8'hC2;
  picture_data[ 7062 ] = 8'h08;
  picture_data[ 7063 ] = 8'hE2;
  picture_data[ 7064 ] = 8'h08;
  picture_data[ 7065 ] = 8'hA1;
  picture_data[ 7066 ] = 8'h10;
  picture_data[ 7067 ] = 8'h80;
  picture_data[ 7068 ] = 8'h10;
  picture_data[ 7069 ] = 8'h80;
  picture_data[ 7070 ] = 8'h31;
  picture_data[ 7071 ] = 8'h63;
  picture_data[ 7072 ] = 8'h10;
  picture_data[ 7073 ] = 8'h40;
  picture_data[ 7074 ] = 8'h29;
  picture_data[ 7075 ] = 8'h22;
  picture_data[ 7076 ] = 8'h31;
  picture_data[ 7077 ] = 8'h83;
  picture_data[ 7078 ] = 8'h20;
  picture_data[ 7079 ] = 8'hC0;
  picture_data[ 7080 ] = 8'h39;
  picture_data[ 7081 ] = 8'h42;
  picture_data[ 7082 ] = 8'h41;
  picture_data[ 7083 ] = 8'h42;
  picture_data[ 7084 ] = 8'h49;
  picture_data[ 7085 ] = 8'h41;
  picture_data[ 7086 ] = 8'h51;
  picture_data[ 7087 ] = 8'h61;
  picture_data[ 7088 ] = 8'h51;
  picture_data[ 7089 ] = 8'h40;
  picture_data[ 7090 ] = 8'h51;
  picture_data[ 7091 ] = 8'hA2;
  picture_data[ 7092 ] = 8'h51;
  picture_data[ 7093 ] = 8'hA2;
  picture_data[ 7094 ] = 8'h49;
  picture_data[ 7095 ] = 8'hA2;
  picture_data[ 7096 ] = 8'h39;
  picture_data[ 7097 ] = 8'h21;
  picture_data[ 7098 ] = 8'h41;
  picture_data[ 7099 ] = 8'h83;
  picture_data[ 7100 ] = 8'h41;
  picture_data[ 7101 ] = 8'hC4;
  picture_data[ 7102 ] = 8'h39;
  picture_data[ 7103 ] = 8'hA4;
  picture_data[ 7104 ] = 8'h31;
  picture_data[ 7105 ] = 8'h43;
  picture_data[ 7106 ] = 8'h42;
  picture_data[ 7107 ] = 8'h05;
  picture_data[ 7108 ] = 8'h39;
  picture_data[ 7109 ] = 8'hA4;
  picture_data[ 7110 ] = 8'h20;
  picture_data[ 7111 ] = 8'hE1;
  picture_data[ 7112 ] = 8'h52;
  picture_data[ 7113 ] = 8'h47;
  picture_data[ 7114 ] = 8'h20;
  picture_data[ 7115 ] = 8'hC1;
  picture_data[ 7116 ] = 8'h29;
  picture_data[ 7117 ] = 8'h02;
  picture_data[ 7118 ] = 8'h20;
  picture_data[ 7119 ] = 8'hC1;
  picture_data[ 7120 ] = 8'h18;
  picture_data[ 7121 ] = 8'h80;
  picture_data[ 7122 ] = 8'h20;
  picture_data[ 7123 ] = 8'hE2;
  picture_data[ 7124 ] = 8'h18;
  picture_data[ 7125 ] = 8'h81;
  picture_data[ 7126 ] = 8'h18;
  picture_data[ 7127 ] = 8'h81;
  picture_data[ 7128 ] = 8'h18;
  picture_data[ 7129 ] = 8'hC2;
  picture_data[ 7130 ] = 8'h10;
  picture_data[ 7131 ] = 8'h80;
  picture_data[ 7132 ] = 8'h10;
  picture_data[ 7133 ] = 8'h80;
  picture_data[ 7134 ] = 8'h21;
  picture_data[ 7135 ] = 8'h22;
  picture_data[ 7136 ] = 8'h19;
  picture_data[ 7137 ] = 8'h01;
  picture_data[ 7138 ] = 8'h21;
  picture_data[ 7139 ] = 8'h22;
  picture_data[ 7140 ] = 8'h21;
  picture_data[ 7141 ] = 8'h21;
  picture_data[ 7142 ] = 8'h10;
  picture_data[ 7143 ] = 8'hA4;
  picture_data[ 7144 ] = 8'h10;
  picture_data[ 7145 ] = 8'hC4;
  picture_data[ 7146 ] = 8'h19;
  picture_data[ 7147 ] = 8'h66;
  picture_data[ 7148 ] = 8'h29;
  picture_data[ 7149 ] = 8'hC7;
  picture_data[ 7150 ] = 8'h19;
  picture_data[ 7151 ] = 8'h46;
  picture_data[ 7152 ] = 8'h21;
  picture_data[ 7153 ] = 8'h68;
  picture_data[ 7154 ] = 8'h21;
  picture_data[ 7155 ] = 8'h4A;
  picture_data[ 7156 ] = 8'h19;
  picture_data[ 7157 ] = 8'h0A;
  picture_data[ 7158 ] = 8'h10;
  picture_data[ 7159 ] = 8'hA7;
  picture_data[ 7160 ] = 8'h10;
  picture_data[ 7161 ] = 8'hC7;
  picture_data[ 7162 ] = 8'h18;
  picture_data[ 7163 ] = 8'hE6;
  picture_data[ 7164 ] = 8'h08;
  picture_data[ 7165 ] = 8'h84;
  picture_data[ 7166 ] = 8'h10;
  picture_data[ 7167 ] = 8'hE4;
  picture_data[ 7168 ] = 8'h10;
  picture_data[ 7169 ] = 8'hE3;
  picture_data[ 7170 ] = 8'h11;
  picture_data[ 7171 ] = 8'h04;
  picture_data[ 7172 ] = 8'h10;
  picture_data[ 7173 ] = 8'hC3;
  picture_data[ 7174 ] = 8'h10;
  picture_data[ 7175 ] = 8'hC3;
  picture_data[ 7176 ] = 8'h08;
  picture_data[ 7177 ] = 8'h61;
  picture_data[ 7178 ] = 8'h00;
  picture_data[ 7179 ] = 8'h41;
  picture_data[ 7180 ] = 8'h08;
  picture_data[ 7181 ] = 8'h41;
  picture_data[ 7182 ] = 8'h08;
  picture_data[ 7183 ] = 8'h41;
  picture_data[ 7184 ] = 8'h00;
  picture_data[ 7185 ] = 8'h41;
  picture_data[ 7186 ] = 8'h00;
  picture_data[ 7187 ] = 8'h20;
  picture_data[ 7188 ] = 8'h00;
  picture_data[ 7189 ] = 8'h20;
  picture_data[ 7190 ] = 8'h08;
  picture_data[ 7191 ] = 8'h61;
  picture_data[ 7192 ] = 8'h10;
  picture_data[ 7193 ] = 8'hA2;
  picture_data[ 7194 ] = 8'h10;
  picture_data[ 7195 ] = 8'hA2;
  picture_data[ 7196 ] = 8'h10;
  picture_data[ 7197 ] = 8'hC2;
  picture_data[ 7198 ] = 8'h19;
  picture_data[ 7199 ] = 8'h03;
  picture_data[ 7200 ] = 8'h19;
  picture_data[ 7201 ] = 8'h03;
  picture_data[ 7202 ] = 8'h10;
  picture_data[ 7203 ] = 8'hC2;
  picture_data[ 7204 ] = 8'h08;
  picture_data[ 7205 ] = 8'h60;
  picture_data[ 7206 ] = 8'h08;
  picture_data[ 7207 ] = 8'h40;
  picture_data[ 7208 ] = 8'h18;
  picture_data[ 7209 ] = 8'hC2;
  picture_data[ 7210 ] = 8'h10;
  picture_data[ 7211 ] = 8'hC2;
  picture_data[ 7212 ] = 8'h08;
  picture_data[ 7213 ] = 8'hC2;
  picture_data[ 7214 ] = 8'h10;
  picture_data[ 7215 ] = 8'hE2;
  picture_data[ 7216 ] = 8'h10;
  picture_data[ 7217 ] = 8'hC1;
  picture_data[ 7218 ] = 8'h18;
  picture_data[ 7219 ] = 8'hC1;
  picture_data[ 7220 ] = 8'h18;
  picture_data[ 7221 ] = 8'hA0;
  picture_data[ 7222 ] = 8'h29;
  picture_data[ 7223 ] = 8'h22;
  picture_data[ 7224 ] = 8'h31;
  picture_data[ 7225 ] = 8'h63;
  picture_data[ 7226 ] = 8'h18;
  picture_data[ 7227 ] = 8'h80;
  picture_data[ 7228 ] = 8'h4A;
  picture_data[ 7229 ] = 8'h05;
  picture_data[ 7230 ] = 8'h41;
  picture_data[ 7231 ] = 8'hE4;
  picture_data[ 7232 ] = 8'h30;
  picture_data[ 7233 ] = 8'hC0;
  picture_data[ 7234 ] = 8'h59;
  picture_data[ 7235 ] = 8'hA2;
  picture_data[ 7236 ] = 8'h59;
  picture_data[ 7237 ] = 8'h81;
  picture_data[ 7238 ] = 8'hAB;
  picture_data[ 7239 ] = 8'hEA;
  picture_data[ 7240 ] = 8'hA3;
  picture_data[ 7241 ] = 8'hA9;
  picture_data[ 7242 ] = 8'h61;
  picture_data[ 7243 ] = 8'hA1;
  picture_data[ 7244 ] = 8'h51;
  picture_data[ 7245 ] = 8'h00;
  picture_data[ 7246 ] = 8'h38;
  picture_data[ 7247 ] = 8'h60;
  picture_data[ 7248 ] = 8'h51;
  picture_data[ 7249 ] = 8'h63;
  picture_data[ 7250 ] = 8'h49;
  picture_data[ 7251 ] = 8'h83;
  picture_data[ 7252 ] = 8'h39;
  picture_data[ 7253 ] = 8'h63;
  picture_data[ 7254 ] = 8'h39;
  picture_data[ 7255 ] = 8'h83;
  picture_data[ 7256 ] = 8'h29;
  picture_data[ 7257 ] = 8'h02;
  picture_data[ 7258 ] = 8'h31;
  picture_data[ 7259 ] = 8'h64;
  picture_data[ 7260 ] = 8'h29;
  picture_data[ 7261 ] = 8'h02;
  picture_data[ 7262 ] = 8'h20;
  picture_data[ 7263 ] = 8'hC1;
  picture_data[ 7264 ] = 8'h18;
  picture_data[ 7265 ] = 8'hA1;
  picture_data[ 7266 ] = 8'h20;
  picture_data[ 7267 ] = 8'hE2;
  picture_data[ 7268 ] = 8'h10;
  picture_data[ 7269 ] = 8'h40;
  picture_data[ 7270 ] = 8'h20;
  picture_data[ 7271 ] = 8'hA1;
  picture_data[ 7272 ] = 8'h28;
  picture_data[ 7273 ] = 8'hC2;
  picture_data[ 7274 ] = 8'h18;
  picture_data[ 7275 ] = 8'h81;
  picture_data[ 7276 ] = 8'h10;
  picture_data[ 7277 ] = 8'h20;
  picture_data[ 7278 ] = 8'h10;
  picture_data[ 7279 ] = 8'h61;
  picture_data[ 7280 ] = 8'h18;
  picture_data[ 7281 ] = 8'hA1;
  picture_data[ 7282 ] = 8'h18;
  picture_data[ 7283 ] = 8'hA1;
  picture_data[ 7284 ] = 8'h18;
  picture_data[ 7285 ] = 8'hC1;
  picture_data[ 7286 ] = 8'h20;
  picture_data[ 7287 ] = 8'hE2;
  picture_data[ 7288 ] = 8'h18;
  picture_data[ 7289 ] = 8'hC1;
  picture_data[ 7290 ] = 8'h18;
  picture_data[ 7291 ] = 8'hE1;
  picture_data[ 7292 ] = 8'h18;
  picture_data[ 7293 ] = 8'hE1;
  picture_data[ 7294 ] = 8'h10;
  picture_data[ 7295 ] = 8'hC4;
  picture_data[ 7296 ] = 8'h08;
  picture_data[ 7297 ] = 8'h83;
  picture_data[ 7298 ] = 8'h08;
  picture_data[ 7299 ] = 8'h82;
  picture_data[ 7300 ] = 8'h08;
  picture_data[ 7301 ] = 8'hA2;
  picture_data[ 7302 ] = 8'h19;
  picture_data[ 7303 ] = 8'h45;
  picture_data[ 7304 ] = 8'h21;
  picture_data[ 7305 ] = 8'h46;
  picture_data[ 7306 ] = 8'h21;
  picture_data[ 7307 ] = 8'h48;
  picture_data[ 7308 ] = 8'h29;
  picture_data[ 7309 ] = 8'h89;
  picture_data[ 7310 ] = 8'h11;
  picture_data[ 7311 ] = 8'h07;
  picture_data[ 7312 ] = 8'h11;
  picture_data[ 7313 ] = 8'h06;
  picture_data[ 7314 ] = 8'h19;
  picture_data[ 7315 ] = 8'h26;
  picture_data[ 7316 ] = 8'h11;
  picture_data[ 7317 ] = 8'h05;
  picture_data[ 7318 ] = 8'h11;
  picture_data[ 7319 ] = 8'h24;
  picture_data[ 7320 ] = 8'h11;
  picture_data[ 7321 ] = 8'h03;
  picture_data[ 7322 ] = 8'h11;
  picture_data[ 7323 ] = 8'h03;
  picture_data[ 7324 ] = 8'h08;
  picture_data[ 7325 ] = 8'hC2;
  picture_data[ 7326 ] = 8'h10;
  picture_data[ 7327 ] = 8'hC2;
  picture_data[ 7328 ] = 8'h08;
  picture_data[ 7329 ] = 8'h82;
  picture_data[ 7330 ] = 8'h08;
  picture_data[ 7331 ] = 8'h61;
  picture_data[ 7332 ] = 8'h08;
  picture_data[ 7333 ] = 8'h61;
  picture_data[ 7334 ] = 8'h00;
  picture_data[ 7335 ] = 8'h41;
  picture_data[ 7336 ] = 8'h08;
  picture_data[ 7337 ] = 8'h82;
  picture_data[ 7338 ] = 8'h08;
  picture_data[ 7339 ] = 8'h61;
  picture_data[ 7340 ] = 8'h00;
  picture_data[ 7341 ] = 8'h41;
  picture_data[ 7342 ] = 8'h08;
  picture_data[ 7343 ] = 8'h81;
  picture_data[ 7344 ] = 8'h10;
  picture_data[ 7345 ] = 8'hA2;
  picture_data[ 7346 ] = 8'h10;
  picture_data[ 7347 ] = 8'hA2;
  picture_data[ 7348 ] = 8'h10;
  picture_data[ 7349 ] = 8'hA2;
  picture_data[ 7350 ] = 8'h08;
  picture_data[ 7351 ] = 8'hA1;
  picture_data[ 7352 ] = 8'h10;
  picture_data[ 7353 ] = 8'hC2;
  picture_data[ 7354 ] = 8'h10;
  picture_data[ 7355 ] = 8'hC2;
  picture_data[ 7356 ] = 8'h08;
  picture_data[ 7357 ] = 8'h61;
  picture_data[ 7358 ] = 8'h08;
  picture_data[ 7359 ] = 8'h40;
  picture_data[ 7360 ] = 8'h10;
  picture_data[ 7361 ] = 8'hA1;
  picture_data[ 7362 ] = 8'h10;
  picture_data[ 7363 ] = 8'hC2;
  picture_data[ 7364 ] = 8'h19;
  picture_data[ 7365 ] = 8'h03;
  picture_data[ 7366 ] = 8'h19;
  picture_data[ 7367 ] = 8'h23;
  picture_data[ 7368 ] = 8'h19;
  picture_data[ 7369 ] = 8'h02;
  picture_data[ 7370 ] = 8'h20;
  picture_data[ 7371 ] = 8'hE2;
  picture_data[ 7372 ] = 8'h20;
  picture_data[ 7373 ] = 8'hE2;
  picture_data[ 7374 ] = 8'h21;
  picture_data[ 7375 ] = 8'h01;
  picture_data[ 7376 ] = 8'h39;
  picture_data[ 7377 ] = 8'hC4;
  picture_data[ 7378 ] = 8'h39;
  picture_data[ 7379 ] = 8'h84;
  picture_data[ 7380 ] = 8'h20;
  picture_data[ 7381 ] = 8'hE1;
  picture_data[ 7382 ] = 8'h41;
  picture_data[ 7383 ] = 8'hC4;
  picture_data[ 7384 ] = 8'h59;
  picture_data[ 7385 ] = 8'hE4;
  picture_data[ 7386 ] = 8'h59;
  picture_data[ 7387 ] = 8'h40;
  picture_data[ 7388 ] = 8'h9B;
  picture_data[ 7389 ] = 8'h05;
  picture_data[ 7390 ] = 8'hEE;
  picture_data[ 7391 ] = 8'h10;
  picture_data[ 7392 ] = 8'hFE;
  picture_data[ 7393 ] = 8'hD3;
  picture_data[ 7394 ] = 8'hAB;
  picture_data[ 7395 ] = 8'h47;
  picture_data[ 7396 ] = 8'h58;
  picture_data[ 7397 ] = 8'h80;
  picture_data[ 7398 ] = 8'h60;
  picture_data[ 7399 ] = 8'hC2;
  picture_data[ 7400 ] = 8'h59;
  picture_data[ 7401 ] = 8'h04;
  picture_data[ 7402 ] = 8'h49;
  picture_data[ 7403 ] = 8'h03;
  picture_data[ 7404 ] = 8'h28;
  picture_data[ 7405 ] = 8'hA1;
  picture_data[ 7406 ] = 8'h31;
  picture_data[ 7407 ] = 8'h02;
  picture_data[ 7408 ] = 8'h20;
  picture_data[ 7409 ] = 8'hC1;
  picture_data[ 7410 ] = 8'h20;
  picture_data[ 7411 ] = 8'h81;
  picture_data[ 7412 ] = 8'h18;
  picture_data[ 7413 ] = 8'h61;
  picture_data[ 7414 ] = 8'h10;
  picture_data[ 7415 ] = 8'h40;
  picture_data[ 7416 ] = 8'h10;
  picture_data[ 7417 ] = 8'h40;
  picture_data[ 7418 ] = 8'h10;
  picture_data[ 7419 ] = 8'h20;
  picture_data[ 7420 ] = 8'h18;
  picture_data[ 7421 ] = 8'h60;
  picture_data[ 7422 ] = 8'h18;
  picture_data[ 7423 ] = 8'h61;
  picture_data[ 7424 ] = 8'h18;
  picture_data[ 7425 ] = 8'h81;
  picture_data[ 7426 ] = 8'h18;
  picture_data[ 7427 ] = 8'h81;
  picture_data[ 7428 ] = 8'h18;
  picture_data[ 7429 ] = 8'h81;
  picture_data[ 7430 ] = 8'h18;
  picture_data[ 7431 ] = 8'hA1;
  picture_data[ 7432 ] = 8'h18;
  picture_data[ 7433 ] = 8'hA1;
  picture_data[ 7434 ] = 8'h18;
  picture_data[ 7435 ] = 8'hA1;
  picture_data[ 7436 ] = 8'h18;
  picture_data[ 7437 ] = 8'hC1;
  picture_data[ 7438 ] = 8'h10;
  picture_data[ 7439 ] = 8'hA1;
  picture_data[ 7440 ] = 8'h18;
  picture_data[ 7441 ] = 8'hC1;
  picture_data[ 7442 ] = 8'h18;
  picture_data[ 7443 ] = 8'hC1;
  picture_data[ 7444 ] = 8'h21;
  picture_data[ 7445 ] = 8'h02;
  picture_data[ 7446 ] = 8'h08;
  picture_data[ 7447 ] = 8'h83;
  picture_data[ 7448 ] = 8'h00;
  picture_data[ 7449 ] = 8'h62;
  picture_data[ 7450 ] = 8'h00;
  picture_data[ 7451 ] = 8'h82;
  picture_data[ 7452 ] = 8'h00;
  picture_data[ 7453 ] = 8'h61;
  picture_data[ 7454 ] = 8'h10;
  picture_data[ 7455 ] = 8'hC3;
  picture_data[ 7456 ] = 8'h10;
  picture_data[ 7457 ] = 8'hC3;
  picture_data[ 7458 ] = 8'h19;
  picture_data[ 7459 ] = 8'h05;
  picture_data[ 7460 ] = 8'h21;
  picture_data[ 7461 ] = 8'h67;
  picture_data[ 7462 ] = 8'h10;
  picture_data[ 7463 ] = 8'hE5;
  picture_data[ 7464 ] = 8'h11;
  picture_data[ 7465 ] = 8'h05;
  picture_data[ 7466 ] = 8'h11;
  picture_data[ 7467 ] = 8'h25;
  picture_data[ 7468 ] = 8'h11;
  picture_data[ 7469 ] = 8'h04;
  picture_data[ 7470 ] = 8'h11;
  picture_data[ 7471 ] = 8'h03;
  picture_data[ 7472 ] = 8'h08;
  picture_data[ 7473 ] = 8'hE2;
  picture_data[ 7474 ] = 8'h10;
  picture_data[ 7475 ] = 8'hE2;
  picture_data[ 7476 ] = 8'h08;
  picture_data[ 7477 ] = 8'hA1;
  picture_data[ 7478 ] = 8'h10;
  picture_data[ 7479 ] = 8'hE3;
  picture_data[ 7480 ] = 8'h08;
  picture_data[ 7481 ] = 8'hA2;
  picture_data[ 7482 ] = 8'h08;
  picture_data[ 7483 ] = 8'h81;
  picture_data[ 7484 ] = 8'h08;
  picture_data[ 7485 ] = 8'h81;
  picture_data[ 7486 ] = 8'h08;
  picture_data[ 7487 ] = 8'h81;
  picture_data[ 7488 ] = 8'h10;
  picture_data[ 7489 ] = 8'hA2;
  picture_data[ 7490 ] = 8'h08;
  picture_data[ 7491 ] = 8'h61;
  picture_data[ 7492 ] = 8'h08;
  picture_data[ 7493 ] = 8'h61;
  picture_data[ 7494 ] = 8'h00;
  picture_data[ 7495 ] = 8'h40;
  picture_data[ 7496 ] = 8'h08;
  picture_data[ 7497 ] = 8'h61;
  picture_data[ 7498 ] = 8'h08;
  picture_data[ 7499 ] = 8'h81;
  picture_data[ 7500 ] = 8'h10;
  picture_data[ 7501 ] = 8'hC2;
  picture_data[ 7502 ] = 8'h10;
  picture_data[ 7503 ] = 8'hA1;
  picture_data[ 7504 ] = 8'h10;
  picture_data[ 7505 ] = 8'hA2;
  picture_data[ 7506 ] = 8'h10;
  picture_data[ 7507 ] = 8'hC2;
  picture_data[ 7508 ] = 8'h10;
  picture_data[ 7509 ] = 8'hA1;
  picture_data[ 7510 ] = 8'h08;
  picture_data[ 7511 ] = 8'h81;
  picture_data[ 7512 ] = 8'h10;
  picture_data[ 7513 ] = 8'hA1;
  picture_data[ 7514 ] = 8'h10;
  picture_data[ 7515 ] = 8'hA1;
  picture_data[ 7516 ] = 8'h18;
  picture_data[ 7517 ] = 8'hE3;
  picture_data[ 7518 ] = 8'h21;
  picture_data[ 7519 ] = 8'h23;
  picture_data[ 7520 ] = 8'h21;
  picture_data[ 7521 ] = 8'h22;
  picture_data[ 7522 ] = 8'h20;
  picture_data[ 7523 ] = 8'hE2;
  picture_data[ 7524 ] = 8'h18;
  picture_data[ 7525 ] = 8'hC1;
  picture_data[ 7526 ] = 8'h21;
  picture_data[ 7527 ] = 8'h22;
  picture_data[ 7528 ] = 8'h29;
  picture_data[ 7529 ] = 8'h63;
  picture_data[ 7530 ] = 8'h39;
  picture_data[ 7531 ] = 8'h84;
  picture_data[ 7532 ] = 8'h20;
  picture_data[ 7533 ] = 8'hC1;
  picture_data[ 7534 ] = 8'h20;
  picture_data[ 7535 ] = 8'h80;
  picture_data[ 7536 ] = 8'h51;
  picture_data[ 7537 ] = 8'h82;
  picture_data[ 7538 ] = 8'h71;
  picture_data[ 7539 ] = 8'hA1;
  picture_data[ 7540 ] = 8'hC3;
  picture_data[ 7541 ] = 8'hE8;
  picture_data[ 7542 ] = 8'hFE;
  picture_data[ 7543 ] = 8'h50;
  picture_data[ 7544 ] = 8'hFE;
  picture_data[ 7545 ] = 8'h50;
  picture_data[ 7546 ] = 8'hDC;
  picture_data[ 7547 ] = 8'h6B;
  picture_data[ 7548 ] = 8'hAA;
  picture_data[ 7549 ] = 8'h86;
  picture_data[ 7550 ] = 8'hA2;
  picture_data[ 7551 ] = 8'h69;
  picture_data[ 7552 ] = 8'h60;
  picture_data[ 7553 ] = 8'hE4;
  picture_data[ 7554 ] = 8'h51;
  picture_data[ 7555 ] = 8'h04;
  picture_data[ 7556 ] = 8'h20;
  picture_data[ 7557 ] = 8'h40;
  picture_data[ 7558 ] = 8'h28;
  picture_data[ 7559 ] = 8'hA1;
  picture_data[ 7560 ] = 8'h20;
  picture_data[ 7561 ] = 8'h60;
  picture_data[ 7562 ] = 8'h18;
  picture_data[ 7563 ] = 8'h61;
  picture_data[ 7564 ] = 8'h18;
  picture_data[ 7565 ] = 8'h41;
  picture_data[ 7566 ] = 8'h10;
  picture_data[ 7567 ] = 8'h41;
  picture_data[ 7568 ] = 8'h10;
  picture_data[ 7569 ] = 8'h41;
  picture_data[ 7570 ] = 8'h18;
  picture_data[ 7571 ] = 8'h41;
  picture_data[ 7572 ] = 8'h20;
  picture_data[ 7573 ] = 8'h61;
  picture_data[ 7574 ] = 8'h20;
  picture_data[ 7575 ] = 8'hA2;
  picture_data[ 7576 ] = 8'h20;
  picture_data[ 7577 ] = 8'hA1;
  picture_data[ 7578 ] = 8'h18;
  picture_data[ 7579 ] = 8'hA1;
  picture_data[ 7580 ] = 8'h18;
  picture_data[ 7581 ] = 8'h81;
  picture_data[ 7582 ] = 8'h18;
  picture_data[ 7583 ] = 8'hA1;
  picture_data[ 7584 ] = 8'h18;
  picture_data[ 7585 ] = 8'hC1;
  picture_data[ 7586 ] = 8'h18;
  picture_data[ 7587 ] = 8'hC1;
  picture_data[ 7588 ] = 8'h18;
  picture_data[ 7589 ] = 8'hE2;
  picture_data[ 7590 ] = 8'h10;
  picture_data[ 7591 ] = 8'h80;
  picture_data[ 7592 ] = 8'h10;
  picture_data[ 7593 ] = 8'hA1;
  picture_data[ 7594 ] = 8'h10;
  picture_data[ 7595 ] = 8'hA1;
  picture_data[ 7596 ] = 8'h21;
  picture_data[ 7597 ] = 8'h02;
  picture_data[ 7598 ] = 8'h00;
  picture_data[ 7599 ] = 8'h00;


  pic_pointer = 13'd0;   
 end                     
 

 always@(posedge CLK)    
 begin                   
                         
  scl <= ~scl;           
                         
 end                     
                         
 always@(posedge CLK)    
 begin                   
                         
  case(state)            
                         
   init:                 
   begin                 
                         
    rst <= 1'b1;         
    dc <= 1'b0;//initialize to low
    mosi <= 1'b0;//initialize to low
    cs <= 1'b1;          
    state <= actRst;     
    delay <= 16'd0;      
                         
   end                   
                         
   actRst:               
   begin                 
                         
    rst <= 1'b0;         
    state <= drst;       
                         
   end                   
                         
   drst:                 
   begin                 
                         
    if(delay <= actRst_d)
    begin                
     delay <= delay + 16'd1; 
    end                  
    else                 
    begin                
     rst <= 1'b1;        
     delay <= 16'd0;     
     state <= ddrst;     
    end                  
                         
   end                   
                         
   ddrst:                
   begin                 
                         
    if(delay <= dactRst_d)
    begin                
     delay <= delay + 16'd1;
    end                  
    else                 
    begin                
     delay <= 16'd0;     
     state <= lc;        
    end                  
                         
   end                   
                         
   lc:                   
   begin                 
                         
    if(cmd[cmd_counter] == 8'h00)
    begin                
     state <= lc;        
    end                  
    else                 
    begin                
     case(cmd[cmd_counter])
      SLPOUT  : params_left <= 14'h00;
      FRMCTR1 : params_left <= 14'h03;
      FRMCTR2 : params_left <= 14'h03;
      FRMCTR3 : params_left <= 14'h06;
      INVCTR  : params_left <= 14'h01;
      PWCTR1  : params_left <= 14'h03;
      PWCTR2  : params_left <= 14'h01;
      PWCTR3  : params_left <= 14'h02;
      PWCTR4  : params_left <= 14'h02;
      PWCTR5  : params_left <= 14'h02;
      VMCTR1  : params_left <= 14'h01;
      GMCTRP1 : params_left <= 14'h10;
      GMCTRN1 : params_left <= 14'h10;
      PWCTR6  : params_left <= 14'h01;
      COLMOD  : params_left <= 14'h01;
      MADCTL  : params_left <= 14'h01;
      INVON   : params_left <= 14'h00;
      DISPON  : params_left <= 14'h00;
      CASET   : params_left <= 14'h04;
      RASET   : params_left <= 14'h04;
      RAMWR   : params_left <= 14'd3800; // Modified for number of pixels
      default : params_left <= 14'h00;
     endcase             
     data <= cmd[cmd_counter];
     cmd_counter <= cmd_counter + 5'b1;
     state <= ldc;       
    end                  
                         
   end                   
                         
   dpcmd: begin          
                         
    if(delay < pcmd)     
    begin                
     delay <= delay + 16'd1;
    end                  
    else                 
    begin
     state <= lc;
     delay <= 16'd0;
    end

   end

   dmw_c: begin

    if(delay < mw_c)
    begin
     delay <= delay + 16'd1;
    end
    else
    begin
     state <= rdc; // Raise dc for params
     delay <= 16'd0; // Reset delay
    end

   end

   ldc: 
   begin

    dc <= 1'b0;
    state <= sm;

   end

   sm: 
   begin

    if(dc == 1'b1 && cmd[cmd_counter-5'd1] == RAMWR)
    begin
     if(pixel_bit_counter == 4'b1111)
     begin
      state <= lcs;
     end
     else if(pixel_bit_counter == 4'b0000)
     begin
      state <= slb;
      pixel_bit_counter <= 4'b1111;
     end
     else
     begin
      state <= send;
     end

     mosi <= pixel_data[pixel_bit_counter];
     pixel_bit_counter <= pixel_bit_counter - 4'b0001;
    end
    else
    begin
     if(bit_counter == 3'b111)
     begin
      state <= lcs;
     end
     else if(bit_counter == 3'b000)
     begin
      state <= slb;
      bit_counter <= 3'b111;
     end
     else
     begin
      state <= send;
     end

     mosi <= data[bit_counter];
     bit_counter <= bit_counter - 3'b001;
    end
 
   end

   lcs: 
   begin

    if(scl == 1'b1)
    begin
     cs <= 1'b0;
     state <= send;
    end
    else
    begin
     state <= lcs;
    end

   end

   send: 
   begin

    if(scl == 1'b1)
    begin
     state <= sm;
    end
    else
    begin
     state <= send;
    end

   end

   slb: 
   begin

    if(scl == 1'b1)
    begin
     state <= rcs;
    end
    else
    begin
     state <= slb;
    end

   end

   rcs: 
   begin
   
    cs <= 1'b1;
    if(dc == 1'b0)
    begin
     if(cmd_counter == 5'd20)
     begin
      state <= dmw_p; // short
     end
     else if(cmd_counter == 5'd23)
     begin
      state <= dmw_c; // long
     end
     else
     begin
      if(cmd[cmd_counter-5'd1] == FRMCTR3)
      begin
       state <= dfrmctr3_c;
      end
      else if(cmd[cmd_counter-5'd1] == GMCTRP1 ||
          cmd[cmd_counter-5'd1] == GMCTRN1)
      begin
       state <= dgmctr_c;
      end
      else if(cmd[cmd_counter-5'd1] == CASET ||
	  cmd[cmd_counter-5'd1] == RASET)
      begin
       state <= dcr_c;
      end
      else if(cmd[cmd_counter-5'd1] == SLPOUT)
      begin
       state <= dsleep;
      end
      else
      begin
       state <= rdc;
      end
     end
    end
    else
    begin
     if(cmd_counter == 5'd23)
     begin
      state <= dmw_p; // Provide 6us delay after each parameter
     end
     else
     begin
      if(cmd[cmd_counter-5'd1] == FRMCTR3)
      begin
       state <= dfrmctr3_p;
      end
      else if(cmd[cmd_counter-5'd1] == GMCTRP1 ||
	      cmd[cmd_counter-5'd1] == GMCTRN1)
      begin
       state <= dgmctr_p;
      end
      else if(cmd[cmd_counter-5'd1] == CASET ||
	      cmd[cmd_counter-5'd1] == RASET)
      begin
       state <= dcr_p;
      end
      else
      begin
       state <= lp;
      end
     end
    end
   
   end

   rdc: 
   begin

    dc <= 1'b1;
    state <= lp;

   end

   lp: 
   begin

    if(cmd[cmd_counter-5'd1] == RAMWR)
    begin
     pixel_data[15:8] <= picture_data[pic_pointer];
     pixel_data[7:0] <= picture_data[pic_pointer + 13'd1];
     pic_counter <= pic_counter + 13'd2;
    end
    else
    begin
     data <= params[param_counter];
    end 

    if(params_left == 14'd0)
    begin
     state <= dpcmd;// need to provide delay
    end
    else
    begin
     param_counter <= param_counter + 7'd01;
     params_left <= params_left - 14'd1;
     state <= sm;
    end                                     

   end

   dmw_p: begin
    
    if(delay < mw_p)
    begin
     delay <= delay + 16'd1;
    end
    else
    begin
     if(cmd_counter == 5'd20)
     begin
      state <= rdc;
     end
     else
     begin
      state <= lp;
     end
     delay <= 16'd0;
    end

   end

   dfrmctr3_c: 
   begin

    if(delay < frmctr3)
    begin
     delay <= delay + 16'd1;
    end
    else
    begin
     state <= rdc;
     delay <= 16'd0; 
    end

   end

   dfrmctr3_p:
   begin

    if(delay < frmctr3)
    begin
     delay <= delay + 16'd1;
    end
    else
    begin
     state <= lp;
     delay <= 16'd0;
    end
 
   end

   dgmctr_c:
   begin

    if(delay < gmctr)
    begin
     delay <= delay + 16'd1;
    end
    else
    begin
     state <= rdc;
     delay <= 16'd0;
    end

   end

   dgmctr_p:
   begin

    if(delay < gmctr)
    begin
     delay <= delay + 16'd1;
    end
    else
    begin
     state <= lp;
     delay <= 16'd0;
    end

   end

   dcr_c:
   begin

    if(delay < cr)
    begin
     delay <= delay + 16'd1;
    end
    else
    begin
     state <= rdc;
     delay <= 16'd0;
    end

   end

   dcr_p:
   begin

    if(delay < cr)
    begin
     delay <= delay + 16'd1;
    end
    else
    begin
     state <= lp;
     delay <= 16'd0;
    end

   end

   dsleep:
   begin

    if(delay < sleep)
    begin
     delay <= delay + 16'd1;
    end
    else
    begin
     state <= rdc;
     delay <= 16'd0;
    end

   end

  endcase
 end

 assign RST = rst;
 assign SCL = scl;
 assign DC = dc;
 assign MOSI = mosi;
 assign CS = cs;

endmodule
